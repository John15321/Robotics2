��   T�A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ������DMR_�SHFERR_T�   $�OFFSET �  	��/G�RP:� �$MA��R_DO�NE  $OT_MINUSJ 7 	sPLzd�COUNJ$REYFj�PO{���I$BCKLS�H_SIG�E?ACHMSTj��SPC�
�MOV�n ~ADAPT_�INERJ F�RICCOL_�P,MGRAV8�� HISI�DSPk�HIFkT_7 O ��Nm�MCH� S��ARM_PAR�AO dcAN�Go y2�CL�DE7�CALI�BDn$GE�AR�2� RINYG��<$]_dΗREL3� �1  	��CL|o: � ��AX{  $PS�_�TI���T_IME �J� �_CMD��"FB�VA �&CL_OyV�� FRMZ�$�DEDX�$NA� %�CUR�L�W���T{CK�%�FMSV��M_LIF	��'83:c$�-9_09:_��=��%3d6W� �"�PCgCOM��FB� yM�0�MAL_�#ECI�P:!o"7DTYkR_|"�5�:#�1END�4���o1 l5M̦P PL� W ݀�STA:#TRGQ_M��� KNiFS� uHYsJ� hG�I�JI�JI�D���$�ASS> �S���A�����@�VERSI� �G�  �i~�AIRTUAL�O��AS 1�H� ��� 	 ��\_G_�_k_�_ �_�_�_�_�_�ZP���i�Y�ABo0l�e������J 9������Zyw�>/o�o+oUl�o@�o�o�o�o�k;�Ar*gyd���d�������=L̙���?����@�=�b�t����������Ώ�����(�{ �US�a�K����D  2���ğ֟���@��0�B�T���<�� ~�������Ưد����� �2�D���Pr�( �x����������� Ͽ���>�)�b�Mϰ��qϖϼ��$4 �12\���P��OM��M���PW�O���/N�=��C�f=�D	�C�4��<E>?,�,>��BQ�ʁB0�@ߙϽ�y�d�>��x$Af�r@��{b;U: :��T�X�At�8�ߙ8X���M濎M�-��4Ђ|�f���?�*��c����LN�ԏLS�FX���� ���T���P�������'���%��345?678901G�O� t�x�q���m������� ����D�}���z� H��lZ|���� �.��2 V h����n@� ��/r�U/�� �//�/�/�/�/8/	? ?n/�/N?<?r?`?�? �?�/�?"?4?�?�?O 8O&O\O�?�?�O�?�? �OFO�O�O�O"_xOI_ [_�O_�_|_�_�_�_ �_>_ob_t_�_�_Bo xofo�o�_o�o(o:o �o,<b�o� ��oP����� (�~O���.� ��� ����܏2�D��h�z� H�Əl�Z�|�����ɟ ۟.������2� �V� h��������n�@�¯ ����r���U����� ����������8�	� �n�пN�<�r�`ϖ� ������"�4Ϯπ�� 8�&�\�n�}��ϕ��͎�0hp����9���$PLCL_GR�P 1S��� D�?�  ���;��_� J��n�������� ���%��