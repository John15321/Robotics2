��  	w^�A��*SYST�EM*��V9.1�0185 12�/11/2019� A  �����AAVM_�WRK_T  �� $EXP�OSURE  �$CAMCLB�DAT@ $PS_TRGVT��$X aH]ZgDISfWg�PgRgLENS_CENT_X��YgyORf  � $CMP_G�C_�UTNUM�APRE_MASwT_C� 	��GRV_M{$�NEW��	ST�AT_RUNAR�ES_ER�VTSCP6� aTCb32:dXSM�p&&�#END!�ORGBK!SMp��3!UPD�O�ABS; � P/ �  $P�ARA�  ����AIO_wCNV� l� �RAC�LO�M�OD_TYP@F+IR�HAL�>#�IN_OU�FA�C� gINTER�CEPfBI�I�Z@!LRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CESI0�!H1�!"PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W� @V�R!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2 � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1 �A�UTOB U��0 9DE7VIC4STI�0�A� P@13��`BQd�f"VAL�#ISP�_UNI�#p_D�Ov7IyFR_F �@K%D13�;A�c��C_WA?t�a�zO�FF_@N�DEL�xLF0q�A�qr�?q�p�C?��`�A�E�C#�s�AT�B�tcbMO� �sE' � [M�s���2�REV�BI�LF�!XI� %�R�  � OD�}`j�$NO`M�^�x�/��"u�� ������`��@Dd p{ E RD_Eb�~�$FSSB�&~W`KBD_SE2u�AG� G�2 "_��B�� V�t:5`pׁQC �a_EDu >� � C2�e�`S�p�4%$l ��t$OP�@QB�qy�_OK���0, P_C� y��dh�U ^�`LACI�!�a��� FqCOMM� �0$D��ϑ�@�pX��OR�BIG�ALLOW� �(KD2�2�@VA�R5�d!�AB * ��BL[@S � ,�KJqM�H`S�pZ@M�_O]z���C�Fd X�0GR�@��M�NFL�I���;@UIRE�84�"� SWIT�=$/0_No`S�"C�F_�G� �>0WARNMxp�d��%`LI�V`NS]T� COR-r�FLTR�TRA�T T�`� $A�CCqS�� X�r�$ORI�.&ӧR�T�`_SFg��HUGV0I�p�T��TPA�I��T����HK�� � ��#@a���HDR�B��2�BJ; �C���3�4�5�6��7�8�  ��0��x@�2 @.� TRQ��$%f��4ր����_U����� COc <�� ����Ȩ3�2��L�LECM�-�MULTIV4�"$��A
2;FS�ILDD�
1��z@T_1b ; 4� STY2�b�4�=@�)24��m9eCռ� |9$��.p��6�I`�* �\�TO��E��EXT���ї��B�ў2�2�0D���@��1b.'�B �9�G�Q� �"Q� /%�a��X�%�?s!DԂU� Sҟ�;A�Ɨ�M8�� � CՋO�! L�0a�� �X׻pAβ$JOB�B����  ��IGO�" dӀ������X�-'x���G�ҧ��C��`��b# tӀF̝ �CNG�AiBA � ϑ��!���/1��À �0����R0P/pY�����$
�|���BqF]�
2J]�_)RN��C`J`�e*�J?�D/5C�	�pӧ��@{ UG�ArzO3л!% \�0�RO�6� �IT<�s� NOM_8pn#��c ���TU��@P� � ��&"+P��� ӨP�	ݭ��RAx@n �3�A����
$TF3%#D%3
T��wpU�13��}�%mHrzT1�E���ޣ�#ݤp�%ߢQlYNT�"�� DBGDE�!'D�]�PU���@t����"��AX��"�uwTAI2sBUFۆ82�?!�1( ��P&�V`PI84'mP��'M�(M�)B �&F>�'SIMQS�@ZwKEE3PAT��zЙ8"�"����Cb��)S�0��`JB���ľaDECg:� g5�Ҳ����* �U�CHNS_EMPͲG$G��7�_�<�c;�1_FP)�TC�6S���5�`%��4�} ��V����W��JR����SEGFRAq�O�� #P�T_LIN�KCP�VF�g��`  C$+ ���ckBZ�PBzr��|�@6,` +� ԦE��A�0��Ad0o`�Ar�D���Id1SIZh���	T�FT�C�Z1Y�ARSm��CP@�'�Ic\1@cX�0<@Lp����0�VCRCߥ�sCC���U1@�X�1��2�Mpq�U�1`��X�Q�UDݤأiC k�p��
DK`݀f��RhEVRf �Fha_
	EF�0N�f�Pd1��&h��5�jC}�+��VSCA[��A��fK2�4��-�	<�ׇMARG���"a�F@@���1DcQ�rN�0LEW�-��R��P<��o�l��RɄ.� ����ǯ��� 5ڡR� HANC��$LG5��a��Ӑ��ـF��Ae����0RYr�3
����
��@ �RA��
�AZ��0Q�N`�O��FCT��sp�F��R�0\P0b ADI��O�� +���+���&���5�5Є���S[�g���BMPUD(PY�1��GAESCPjc��W��%N  S-��U0ۑuU�/)�TIT'q�<�b�%ECA:!�!E'RRLd��0�&Q��OR�B$������~�0$RUN_O��SYS��4������u�REV�d@��?DBPXWO�P�=10�$SKo�"�1�DBT�pTRLn�2 �C AC��0��%�m�U DJ�p��_�`�!A�ǀM�P5L�A_2WA��j�EE��D!w�!%R|hO�UMMY9��ڠ�1� ��DBd[��3���!PR�Q? 
�Dٱ9���4 г$�r�$ Q��L�ة5寣�����6��z�PC�7�*�z�PENEC0Tq8I�����RECOR$�9�H m��4$L��5$أ�"E���0R@��VA��_Dց� gROS) �"SK������I�=�א��P�A��JVBETURYN���SMR(�U) v#�CRʰEWMDB=0GNALV �"�$LA� [�*6{$P-�7$Pv�Fs�8o�!�PC��#�DO^@-�Ŵ��|�R˶GO_AW�FܱMOz��p���CSS_CN4�Y�O�:��T��0���I�D�T�2��2�NB��O@�J��v`Iְ� ; P $f>�RB�B��PI�{POl�I_BY���vЅ�TVR��HND=G$�< H�`�1�a�@cS��DSBL�I��s���0}���L�S$�=��0� ��FB�FEձL�9�����5��>D�$cDO�1�C�pMC�0@q��4��9�RH��qW��K4ELE�u�r���SLAVr?xBINS ���#t����_R@P�@ \`�pS�}�l�}�l�{u���[!e��ے�I����B��W��D�N3TV�#�VE�$��SKIlA4;3��	2UB�1J�f�1C�
D�SAF7�5��_S}V6�EXCLU-�:�XrONL�0�YY��s����HI_yVՀ�RPPLYo��RCsH� �0_M��Q�VRFY_�I�.Mms$IOv0��}��1UB���Oj�3LS����%4!��:@��P�$�ĆAUTOCNE �����.��GCHD�s��_ؤ��3s�AF��CPDe�T!��_�G Ao���_�0�  ��NOC�tBxB�pT��A ���z�SG�` �C � 
$CUR8�U��!" �� �T@B�����ANNUNC�#���䱐b���()%!��X-*I&�EF��IC�D @�`F
"a��POTX�aө������ؿ��֠EM��NIBߢE�·"�G� A���$DAY��LOA�D`Ԟ��"��5�����EFF_AXIJ�Fo�%Q�O0|�:�_RTRQV1�G D�a��?0�R�K3�0S45 2Fpz@]w:1a��A0p�/1sAH 0B!�1A0�T�2�ûvDUX��u]��CABsAIs"f�pNS�1�PID�@CPWSs�5�AWpV`��V_�0q0�P�DI�AGysAJ� '1$VX��ET	`�U rT��EJ��{RRf��!��TVE�� SW|AZ�sP�0�:5q0�G}P:1OHP5�1P�P|@�SIR|�{RB �P�2�3%qZQC �B B��H�^��E`��5q0�I��?0���URQDMW�EMSB�?UA�px�EjB�TLIFE�`K#iP��uRN|QFB�U@%!zSFB�a�%"C�+��N��Y'p�gFLA�t& OVڰ�VHE��BSUP�PO(��uRI�_�T��Q_X�d��
 gZjWj� g��%!��6�XZ*�ϡfA+Y2xhC��T�㰢DEN�pBE%!J�� ��F_8p�A���p��K `Q�CACH8�*r�bSIZ�V�P�`�N��UFFI`�oP�ឤ2���6����M;��tL� 81 KEYIMAG �TM��!�^q�:�Yv����OCVsIE�@�qM ��⼠L~��;�?� Q	��р�dNG0��ST��!�r���t����t0�t0�pEMAIL����!�5/FAUL�"O�r��/���COU��쑁��T��)AP< �$9�p�S�0�0IT��BUF�g;��gEԔo�e��PBe�p�C�:���:�|�G�SAV ��r�[@�b��@ˇÐ�)&P��p印�D��_0e���� �OT겮���3Pm ��0�z3�AX�#f x Xe�C��_G|S
��YN_\�A��Q <I0Dk�TO����BM�2�P5T� F�$�DI[E7�����IR��$ G���!&��Ǳ���:�9�Sa����-��C_ᰂ��K�$�����RpVq���DSPnv6�PCe�IM��\���<�3@U9��P�] �IP���A�`�[�TH�`3�O�0T��\�HSȓ>�BSC���`e�V��
���#���*4NV��G ;���`Y�e�F|A}�ad>���Z��SC%B�a��MER)�F�BCMP)�ETn�� TLrFU`�DUY���R�mb�CaDR�ܠ'�"���SNO�n!UG0*А���%���%P���C"�
ō-"2��|:�o VH *
�L��)�9���G �� ��}�Z{ƥ!{�1{�P1{�6q{�7x�8xɡ9x�|PzȄ�1��1���1��1��1��1���1��1��2��2T�ˑ�2��2��2��U2��2��2��2�ʕ3��3��3�˞�3���3��3��3��3���3��4��61EX	T6An!W��߸���V���uş����@F{DR%DXTE��V� .�uR�
�uRR�EM^@F���BOV�M5�*�A3�TRO�V3�DT��S�MX�b�IN3��PR�"AINDq�cB
��ɐ}���Ge��C\�p�UkA9DO6\�RIVW�R��BGEAR5�IObEK#�cDN��1�`X� zp`dCZ_MsCMp`uQ �F�P;UR��Y ,����? �P>?\o {A?oE� Dw��������Z9pj*PPM�2@RI��<pr�ETUP2_� [ 0q�TDʠ�1p�T������1r�BAC��\ QT�pr��)�%w#8@ó�TIFI�A��0��d��@/PT�B�q�FLUI�t] 1�@�x;�UR�A����R�Б
��:C_0I��$�S_?x��J�CO��"�V�RT��� x$SHqO^14 #�ASS�p-��U̠��BG_ � !.�!��!��!�ÏFORC#�U jD�ATA)A^�rFUZ1��]#2��5�iܖ`)A_ |��NA�V=�������S��S$VI�SI��SC=�SQE� ��5V� O�1�&1BF�4@�&�$PO� I�A��FMR2��` ���2��� 6�!3J�)�CE�#�_����_@IT_Yִ]@M�������DGCLF�EDG�DY�8LD���5@�V���T̐0�ua4��v9 T�FS
��tb P��RB��>}�$EX_RAiHBRA1Y�X��RS@3�K�5�F�G&�	5c Y�� ��SW��O0VDEBUG$�A(��GR� opUz�BK�U��O1M� �0POZ0Y�@���E:�@M�LOOM�9QSM�0E��J���P_E d rp^��TERM[UedVN� ORI֑`PfdV?$�SM_��B`PgdU��Q �XhdV�T UP�ri� -���2d�rS�P�e� G�Z @ELT�O���A�FIG��bZ �Agp�T�Tf�$UFR�$`��aM`ѵ�0OTZg�A�TA��lcNSTאPAT��`�bOPTHJ�ϰE�p8�ذbART؀"ep)�؁���REL�j�SHFTӢ�a��h_�R��̳�V �P$�Wph�1�����t�SHI�`�4Uz � ҁAYLO�� m���l� ��a}!�ޠERV��Sq�x ��hgא�b �K�u.��KRC��ASY1M���WJ+g�Ⴃ�E��a�y�ұU��א���e@�v�eP���ppE�2vORאML3G GRJQ
4jX"��B0V�`G`l�u HO�6Dk ��aN� ��OCaQ@$OP�$e�i��#����Հ�RY��aOU��c�PTR�e����a�e$PWR��IM��rR_˃�d� �P̛cUD��cSV����֔l� $�H�!��ADDR
��HMQG�b������p����!1m H��S���! ��.�畞Ì畫�SEz1�#��S<ܰ
3n $� À�_D��P�.�PR�M_�"LOG�_HTTP_��H1wo (��OBJ� l��$��LEyc���d�p � \�睱AB_��T@SⶢS���{KRL~K�HITCOU�  À�!퀶������M�SS��v�J�QUERY_FL�A!a��B_WEBwSOC�"�HW���a1q�7�IN'CPU�B�!Ou�ˡ��Č������������IOLNr �8��R	� $S�L2$INPU�T_PQ$�ܸP��# ���SLA.�1 sðٿ�p��s��r����^C�F_AS8Bt�$_���[�Nq �!]�/a�ɳ�@ҳUp�HY���l� �F�UOP5Eu ` X������ā������P�����������Ə� M�qqv �l�@;sTAkr��A�TI��.�a�Z0Sն�`PSR�BUZ0ID~0��z���y՜Q�!�u�z`w�3��f�G��N��Z0����IRCA��� �x Ĩ��CY�EA{���!���%�R�`�q|�8��DAY_��}�NTVA���i�¦eu��i�SCAepi�CL��������� qy`���ԧb����N_ՀACQ�Ђ�W�rz� O ��������y�G�<]�O! 2yUQ!҄q{P���P�L�ABzan�Z0t�UN�ISb�PITYX��"ѳ����R$�6D|R_UR�L� �$AL10EAN�@�� �PH�T�wT_U��Jt�q} X��"t�R��" �0A�D�2,J�8FLt@��80
K�3
�UJ]R	5~ ���F|@�1w�FgwD��$�J72�O!�$J�8�	7�@\��7�s�� 8�	�APHMI@Q��Df@�J7J8�
L_�KE��  ��K��LM��  <��XRK��� ��WATCH_VA��!pp��FIEL�D��y`�&��� č0paVyp�ֆCT`��E��BD�LG���� !��LG_SIZ���@��3@�O��FD�I ��,Q��]P�� ��J&3@J&O�J&��J&]PJ&�q�E`1_�CM^c�!{@�*h1F ��'�$��(�#r��&3@�&O��&��'I�(�(,P�&�]P�&�RSI�` 7 (�@LN��B�����@{A� g1��K�u1��L~3t27DAU�5EAS������2�0GH����_��BOOܑ��3 Cr�[�IT8��4�<`n�RE(��8SC�R� ڣs�DIm�S�G`G@RGIPR$D�/L�f�քYB��[�S���Z�W7D[��4f�J{GM�GMNCHH�&[�FN�FK�G��ƶIUF�H2p�HFW�D�HHL�ISTP��JV�H�P�H�0�HRES3YHJ��Kc�C4t@S�f�x�kG�YUJ���DjG 3yE�{��BG�I�`PO�WZ&ES̤"�DOC���FEX.b�TUI�EI/ �� �/!�dDa�CNc�@��p�� 4	��EpA;NOGfANA[�ā��AIt瑜��D�CSZ���c���bO��hO�gS?��b�hS�hNHIGN����0�A�(��dDE��pTLL�qC�1��*�i����T�"$����}�����SA������ʰ��Z�� *�P1�u2�u3�q��8�R�`*І ���V��c��5�z�x�6���P�6�.�ST��R�0Y��`Q� �$E_�C_���I��n���� �sG�*Ї Lo���瀖�x������_�ENS�_���pB~C_ � =��h0Y���@��M�Ch2� ���C�LDP��TRQ�LI��D�2�FLAGZ�2�3�f���Du�f�`�LDf�P�f�O�RGjQy��(RESERV��Ŕ��Ŕ��
#�3�� �� 	O�jUA�f�SVHX0D�R	���'�RCLMC5�şןG���'���MՠJ�/��3$DEBUGMAS��S�D�"R��T�`p�E� TZ��G�MFRQ��ߌ � �HR/S_RU��ځ�yA)��UFREQ� �J�$``�OVEARh����v|P�A7EFI��%���䘡���ѣ� \8 ��$U��g?����PS�p
7 	�C�06�BҒ��G�U�Н�?( �	_1MISCi�� dq1�RQ5	f	TBB@�� ��aa�AX9�!	�"�EXCES���۳)M��.����9���ܲSC� � H���_G���,�P�� �2�q�K���|�أB@��B_�FL�IC��B@QUI[RExSMO��O���d�p�L܀M��� �
��19Э��5���pMND�1e�/��o2f2�x�D�#�4I�NAUT(A�4RSM� ��pNZ�b!�Sz^�d�PSTL.w� 4��LOC��RI1P�EX��ACNG�b����b Aե���p�x MF�%7�+�ۂ�P�8e�c0��SUP��FX/ IGG�1 � ���ۃb!C ۃ�Vۄ��V�P���R� ��R�����SD�w��CTIj���c M n��� t-�MD*��)8��`C�L�@�H8�C�DIA�D�2 W]AC��q��C�D��3)!�Oh�/�[ a�CU�V��(����OPA_��.� �t �7㉠f��
 ��P��>P���P��KE�RR�#�-$B�����ND�2N�ND2_TX�XTRA�cp`�M�9�LO�0/�_�L���G�i2����k�RR2൜O� -��1A$�� d$CALI���c%G�a�2�pRsIN�!�<$R� �SW0S� `�ABC>�D_JV �����7�_J3K
E1#SP���PEl�3k�񱀦��J�`����OiqIM<`�'�CSKPS��H� �c�J�1'�Q��%�%'�_AZ#��=!ELNq�N�OCMP�(���z0cRT��h#�1�����1��(o`�*Z��$SMGMP�%�J�G�SCLB���SPH_�`�+0�#\ z��� RTER���`� _�`��*�AP@G�'�4DI�S!�"23U�DF�o�<1LWB8VE�LD�IN��Z`e0_�BL�`��m4���J`]4r7�7�4� IN� �������5QB���t�1��_̰ ��5 �2#5p��4z�936��DHB�r ����p$V� ���#�oa$� �����$\�ൡH �$BELN |��!_ACCEs1� �H`��@IRCi_0���NT���/�$PSB�7�Lo���DL��0�G3ဿ`�F;�I�G�C�G3�B��E�_�qPB-P3Q�����A_MG��D1DPQ2��FW���`�ClU�C�BaXDE�[�PPABN�GRO� EECR�q�_D�!��q�����Ao�$U�SE_� �cP�C�TR�dY�Pb@"� ��YN߰Aa`f��Z�aM����bJPO8_0�AGdINC�����RpT�ig��ENC0L��A�B��@IN7�I�B�e���$NT]3�5NT2c3_@2���cLOQ0���`-�IP����fF0@����� ���e��C�0�fMOSIUQ�����3Q�'�PERCH#  s+�2 ]w� hs��r%���c'["eH
P2P�A�B�uL�T �����e��z�vvgTRK�%ʁAY� �s��,��B;�0��n&8��wbȠMOM���@�»������S�G���C�R� DU�(RS�_BCKLSH_C�B����<v,�"c���݃�b�1a%CLA�LM�d��m�@�C�HK��NGLRTY��5�d����9_Z�1t_UM��l��C��^Q�!����LMTh_L��V#��j���E��Ð�����E����H}���r��xPC�nq�xH���TUl�C�MCv^PbWCN_b�Nuc��SFtA�yVb�g�!8��Bܧ�<�CATs�SH Z��bT�f]����f�0�A�	� QPPAs�gb_Pr�V�_�� 3�`Qp�C�U�F�JG>��X�I�K0OGV�2TORQU�P�/sL���P��Gr1�P��_W ��,��!QAٴBCصHC�صI�I�IHCF�$�˱�-��ZPVC"�@0����N�1T�RP8h�$!Z�JRKT̙�,�ƴ�DB� M���M��_DLBA�rGRVߴ��BC��HC���H_����@�CO1S�p �LN��6� W�=�B@8ٵ 8�
�tڈb�(���Z1�Gv��M�Y?Ѳ��='���T�HET0uNK2a3HC��<C@�CB�kCB<CC� AS��'�
�5�BC5��SB8BCS��GTS��QCo/��'��'��q�$DUC��w���(t5��5Q�q_��+NE��AKS�z)!8 @��A���'����LPH����e��SW�o�b�o�q��⠀֙�����V@�V�5�2@X�Vg�Vt�V���V��V��V��V��H@�Y�_W�ܡv�t�H��H��H��H���H��O1�O@�OT�	V�Og�Ot�O��UO��O��O��O�ցF��"�~bՃ3�S�PBALANCE�_�ѮLEj�H_��SP�1S��b��>q�PFULC�"��"q��:1�|!U�TO_>�F�T1T2B)�B2N%��B�` b$�!f� ���B}C���T�pO@�AɰIN�SEG�B qREV8�& p�aDIF��9�1��'B1��`O!B�!	��Ó�2���`�0���LCHWAR̬R	bAB%���$MECH+���9a?1T�AX9�P�X6�#B7 � 
Y2��{An�eROBQpCR�rX�5M��0�CyA_A��T � x ?$WEIGH6`�#$1��3X�I6a�`sIF�QjPLAG'b��S'b� 'bBIL�EODo�#p�2STD�@�2P�!	��0
`@(Ơ�1�0��0
�`yB<(aA�  2�.t�6/DEBU�3L�@<B=��MMY9�E� qN��D�$D�A�xq$�@S���  �DO_�@A�1� <�0VFL HU�(a�B&B@N�cR�H_p(`GCBO� �� %��T�`�a��T�!~D�@�TICK�30T1"�@%NS��WPNQp1 �CQpRԀ(a!2iU!2|uU�@PROMP6c�E� $IR���&aL��R�p�RMA�I��aa8b�U_@��S� B�:`R��C�OD[CFU.`�6I�D_ppe� �R�G�_SUFF
� �Ca�QdRDO`lW� mU @lVGRC !2Id�SUd!2`e!2leP��Id�De@��0H� �_FIZA9�cO�RD&A �0�B3�6��b&a�@$Z;DTe �CA�Eߦ4 *�!L_�NAQWPriUDEF_I)xr�V5tuU -BhV7DhVasuUou�VIS�����A��hT�s"uS3t���D4l���B7BD5 ���t[CD���O��BLOCKE �Cci_{_�W�qIbC`UMHerIdasIdou Id�rUbK�TeDsUdt Ub5F���q`c,0B�`e r`eas`c���EhP�P� �t,P�q��@W�*�)� �����TE��D� }ALOMB_C��^�0�2VIS!�I�TY�2AS�O'CA�_FRI2#��� SI�q���RTP��_PR��3tC�2W��W���������_��jaEAS�3jbd������p�R���4��5��6�3ORMULA_I���G	w� h ��N7�ECOEFF_O;Q� ��;Qr��G��3S�0�BCA� �O�CCAGR�� � � $ �4u"�BX+PTM��` �AR(�%��CER� qT	�t�`�  +"�LLkd�pS�_S�V�tw�$L��`����v��`� ��SwETU�sMEA�P�(`F��0CA�b�0� g� ���0 �@�o��Q2��q�rHWP�q��tբܑubÕQ�p�q�p+�t��� �PREC�av�pSK_���� P�11_USER^!�"}�08��}�^!VEL"�}��0��!1I�`J ��MTQCFGs��O  YP� OG2�NORE�0P����0��� 4 pݳB7�2H1XYZ�c�J!o yCH0
��_ERR�1� �I�Q��Pۣ@�aAi�����@BUFINDX������R� H�0CU@�QH1���Q��a���"�a$${0��~q��f�o ���G� � $SIj����P�!���VO����0OBJyE���ADJU�B��� �AY�p5��D.�OU�`Վ�'a�b=��T� ]��\��BDIRa�i�� 8��"�0DYN쒣2��T6 �R��,P&@~��OPWOR��� �,�@SY�SBU �SOP���cҎ���U��� P ����PA����C2�OP^`U�!���!XB�AI�IMA�GS��0U�7BIM���o�IN��@�n�RGOVRD��	��K�PM�m�0� ߀�s��H2L�B=з �PMC_E�`cъAENM��A�B1�B7 ���SL�t��� ��0OVSL:�&S�DEX�q}p"/2G2� ��_��G �`��G�`Qfa�B�C�0p�%�c��/_ZER�����s�� @вb5O&`RI��s0
��P��	�� 	��P�L�Ĵ  $�FREE��E��Q	f��!�Ls����yTD0;@ATUS㰎�AC_T��r�UB �_H��s�A4�`t�� D�AI�2RL��a2S�an S���XEY����1�� �0XUP��p��qPX�PF�D3������PG�Ÿ>��$SUBGb5���G�JMPWA�IT�V_%LOWp�BQ��@CVF�Q�ZPG2b!Rz���U3C�C� R��MR�'IG�NR_PL�DB�TB;@P�qH1BW��P�$��UP�%IG�0�PIG3TNLND�&2R�����N�P�)PEED�8HADOW;@������E7S4F1!4pSP]Ds�� L�0AV�05ps0�3UN�0"+d0!R��LY�`�� Q�P��v1��G�$��M�P�@L\+�NPA�T�2�xD��PIP%w0�>��ARSIZ�T���c|q�Om`�h�A�TT���"\�B$�M�EM�B�A>C�3UX���e�PL`�ļ� $���SWIT�CHZ"�AW��ASr�B�BLLBv1��� $BArZ�D�s�BAM� h���I��@J50�����B6�F�A_KN�OW�3R��U!�A�D�H۠~0D��5YPAYLOA鱱�SS�_s�\W��\WZYSL�A�mpLCL_�� !���R�A����T���VF�YC�K��Z貓T��I�XR�M��W_ҬTB���JL�a_J�Q����AND^�9�8d�R�Q����PL�@AL_ ��@~0���A��k�C"�DXSE!��sJ3M`af� T���PDCK��r�C}OŰ_ALPHqc��cBE��W�qo�l���Т�!�� � ��40R_D_1YZ2�TDŰAR�4x!uxEv0s��TIA4_yu5_y6"�MOM��@ks�sxs�s�s��Bv �ADks�vxs�v�sPUB��R�t�uxs�u��r��Bp��� L$PI�1s���^W.��xY.�I:�IH�IV�<p}Q7��!�� !��b�ӆ��73HIG�C73w%p4 Іp4w%� z�І�߈�!!w%SAMP ���B�ЇC�w%�@>c 5�q���7 �� �� ��p0"p��0p�Ҁ����hp���	���INќ�&�ؘ��ϔw"�ښ���:�GAM�MƕS[%�$G#ET��o��D�d��M
ϡIB��2I0�$HI�_��sЩ���E�м�A��٠ʦLW�����٩�ʦ��b��0caC�%CH�K��� 	��nI_ %�����\bxΑ�����s���v���c {�$�h 1���}I� RCH_D��0'� �$)�LE��������hذ�0MS�WFL�$M�`SC�R
(75_����3 ��dƧ���kp��x�p0��DSVv1�P���v�Kǿ�	���S_�SA�A�����NO�`C���d���� d_v_\�J�:ۂ�+R��w�0sD<�4���40�� zʴ�ʈ��چ�1��� �ՕәS�Ak0L���� � ��YL,�a������-��� -���b��9�az�HK����W�{����py�Ȳ�M� ��P��`a�$ 7��"r�M���� � �$���$W���ANG]�Q���d���d@���d���d� נNPP���C��ϐX�0O�c�ΑZq��� �� -�<�OM��"���1�C�U�g�bpCON���0}C�a_�B� |�a�����y7xs7 �s��dzdO~z�A��� �0����0�PP A�PMO�N_QUG� �{ 8�0QCOU��nǀQTH� HO&�n� HYSD@ES�BF� UE� ��@O5$�  �@P�৥���RUNZY���O��� � POP+�%����2ROGRA(��x@:�2�Ov+�IT�xINFO��� �A_��8���`��� (ʰSLEQ�����0�b�`EDd � '� ���r�K�QI#5��EȠNU'(�AUT��%COPAY�Q��8,���M���NB F+U�PRUTZ� I"NF2U�B�$G0�$��RG�ADJ!�BX_��2$�0�&~��&W�(P�(��&73� z�NH`_CYC��ARGNSD9���LGOb��`�NYQ_FREQ��rW����^1RD)L��P:BV0�!�s���CcRE���c�IFH��jNAK�%�4_}G�STATU <å�MAILI�S�&@V��ǀLASTx�1�a04ELEM:1w� �EaNAB��0EASI&A��v� n�?�B���GF�����I���U2���� L�|BAB�C	PRS�LV	A�Fa�I���q1U����JP'c�F?RMS_TRvCΑ���Ci����A�D ��04��& 	~SB 2�  � V��9V(b8WR��R0NTdW&�
�DO�P�W�}�
�22PR �;0Ҟ�GRID}�B7ARS��TY'C��r��O�p!� E_�4!� �R�TOo�>74� � |� �PORXc�	bS�RV�0)(d fDI��T!pAaTd��^g���^g4\i[�^g6\i7�\i8@a��Fj�:1�~$VALU�C���9D7@�F65��� !"E��l�S�1��_@AN���b�1�R c17ATOTA�LH��qCsPWK3I|�QYtREGENWzlr�X�H@c5v�� TR�C�Wq_S���wlp\CV�!���u���1GRE5C�P�p6B+.  sV_H�P�DA���p�S_Yh�i�o6SV�AR���2� �"IG_CSE�3�p b�5_/��tC_�V$CMP,���DE�M����Ie�Z��^���F��HANC�� p&Q$E�2���GINT?`iq��F%��MASK=��@OVR�P� �P��1�Α�W!;�T� �4� �_XF�{�V�P�SLGV�:1� @�K��p5a���ApJpS8h��4��U>�!̬���TEa��`���`�U�Jd���3IL_M~4���p� TQ� ����@-�*\�V4�CB�P{�4A�L�Mc�V1b�V1�p�2�2p�3�3
p�4�4p����p:�`���p��j�|�IN�VIB��<�)���0�U2,�28�3,�38��4,�48� hR�S���� �T $�MC_F�  �B��L����ׅ7pM8�1I׃���S ( �����n�KEEP_H/NADD��!ﴙ@��C��0��Q��?��O��| ���p��܇�REM'�@�IqbL�c�h�U�4�e�HPWD  ;�SBM��P?COLLAB��ph��5q�2�IT50�`�W"NO��FCAqL��� ,���FL�A$SY�N���M� Cq��~XpUP_DLY!=�DELA?�Jq��2Y� AD��	� QSKIP��� �`-O;�NT�yQi�P_-V�� ^U�*����q���q�� u`�ڂ`�ڏ`�ڜ`��Щ`�ڶ`��9�!�J�2R0� �L�EX�@TX3N�7AN� ��N�}�`RDC���� ���Rz�T#OR� ;��R�1��x���;TRGEA�r8h@��RFLG�^��5�ER���SPC��1UM_N��2/TH2N�Q�A� 1� �E�D�Q62 � D�Kш��@2_PC�3]�S���1_0L10_C}2�`2���7 �� $b�  ���	V=�����0 �� �� Sb����mrj��C 2��=��ID� Gy�XUV�L1a�1n��� 10c�_DS��=��a�P�11!� l������#C��AT E��$�Q��bf���;T�3�HOMQE�,0f2n�t`����� ��
i3n��'L9K 0�i4n��n����� )i5n���@/!/3/E/c�f6n��h/z/�/�/�/�/ +f7n��/�/�	??-???Q78n�b?t?�?�?�?�?W%S|���!�  �A�g�p��3�c�Ed�� TC�tD:vtCIIOꑔII@f�O��_OP�E�C4r��}��� WE�� �^@�l�4t y���B$DSB��GGNA��3s:�C��a/�S232zE� ����5���I�CEUS=sSPE|(��aPARIT ��2qOPB���bFLOWO�TR9@?rt��UX�CUuP���aU�XT��a�ERF�ACZTT�U.p��SCHa� t�఩�_`Py���$L ��pOM8���A��8�𥀯�UPDư��f�qPTU@��EX��8#hc�EFA8������RSP�P�a����`�7$USA����9��EX�PIH��(`�pY�eR_$�0q�`mQ�fWR�O�ID���f��FFR�IEND���0$�UFRAMc�pTwOOLvMYH���rLENGTH_VTE�dI�;s��$Z pJxUFI�NV_^ ��_AR�GI%���ITIĨ�BwX�Sw�vG2�gG1�aꀎc�r�w2�_r�O_XP�� �2+q4���N�Sc���C�Pr�q� �G���Rǁ󐒧�XQ؂���h�U���U�������PUd�X �m`E_MG`CT�cH��h���U�dSc%G�W�`ć��ل	D]и@KȅJӂй�������$-� C2���an �i1�h��`2�k2=�3�k3 �j-����iK���F�`�l��`x�|�NtV�uVD��Pq�,��r�P����V������R� �pr�.���E9�<�8Os)E$A��T�CPRh�U�k�ǓS���P���"Sb;Q�! ! �ႃ"��K�锂"���S`�p�p��
_�$$C��S��O����9�9�� ؠVERSIܧ`���i��I#PP��AoAVM_�a2 �� ?0  �5�V�rb�S��� ��A	������9� �����ζ����ϧ�`�R�d�l�0�BS^ �r1�� <@ϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����|»CC`XLM�@v����  d��IN����qEX$?��2_`=�r ���0�IOCip,q ��PZXQ���{�IO'PV �1=�P $-��`ұ�!̺ �?�� � ��//%/7/I/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�o�o�o�o �o�o�o#5GY k}������ ���1�C�U�g�y� ��������ӏ���	� �-�?�Q�c�u����� ����ϟ����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i��{ύϟϱ���� LA�RMRECOV �I��LM_DG �����_IF ���p߂ߔߦ߀��^���������, 
 �G���@�m�����$_� ������ �2�D�V��h��NGTOL � I 	 A�   ����� PPINFO %� $������  1�I
�8 r\������� &W�p�Rd v��������//*/x�PPLI�CATION ?}����LR Ha�ndlingTo�ol y" 
V�9.10P/25���5'
8834�0z#�*F0�!�/1�31y#�,�/�"7�DF1� 5,y#No�ne5+FRA�5/ 6�-B&_�ACTIVE�� � [#��  X3U_TOMODb0)����U5CHGAPO�NL�? �3OUPLED 1M�� �0�?�?�?O;�CUREQ 1	�M�  TIL�L	XOiE_ ~D�wB�m%�MDH6E�2cJH�TTHKYwO��D\COUO_�O7O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q� c�u�����󏽏Ϗ� ����)�;�M�_�q� �����˟ݟ��� �%�7�I�[�m���� 믵�ǯٯ�����!� 3�E�W�i�{���翱� ÿտ�����/�A� S�e�wω��ϭϿ��� ������+�=�O�a� s߅��ߩ߻������߀��'�9�K�CET�O��d?X2DO_CLEAN�?V4���NM  �� O*�<�N�`�r�NDSPDRYR��&U5HI�0�@��� ��&8J\n�����R8MAX@I ��|�~A�7�X����!�2�!X2PLUG�G�0���3t5PRC*��B������.O3����SEGF�0Kz�������//&/^�LAP����Cz/�/�/ �/�/�/�/�/
??.?�@?R?�3TOTAL���3USENU
��; ��?~B@�RGDISPMM�C��AC��@I@���4O������3_STRING� 1
�;
�kM�0ST:
)A�_ITEM13F  nT=OOaOsO�O�O �O�O�O�O�O__'_�9_K_]_o_�_�_�_�I/O SIG�NAL-ETr�yout Mod�e4EInp�PS�imulated�8AOut�\�OVERR�� =� 1007BIn� cycl�U8A�Prog Abo�rc8A�TSta�tus6C	Hea�rtbeat2GMH Faulug~cAler�i�_�o �o�o�o�o $6H ��/K��AO K������� �)�;�M�_�q�����৏��ˏݏ_WOR �/K���=�O�a� s���������͟ߟ� ��'�9�K�]�o�����PO-Kia��-� ��ܯ� ��$�6�H� Z�l�~�������ƿؿ����� �2ϴ�DEV��]�ЯJτϖϨ� ����������&�8� J�\�n߀ߒߤ߶���>��PALTu}� -���)�;�M�_�q�� �������������%�7�I�[�m���GRI� /K�������� ��'9K]o �����������0Ru}I��# q������� //%/7/I/[/m//�/�/�/7PREG �� a�/?'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OGOYO�]��$ARG_�D ?	����A��  �	$�V	[��H]�G��W�I�@S�BN_CONFIQG�P�K�Q�RQ��ACII_SAVE  �TQS�@�TCELLSET�UP �J%  OME_IO�]��\%MOV_H8VPi_o_REPL�_��JUTOBACK�AQ�IQF�RA:\�+ X�_�&P'`T`�'�h� k
P �18/02�/09 11:0/6:04�&�H�-`{o�o�o�o�\���o�%7I[�&� �o������n ��+�=�O�a�s�� ������͏ߏ�|���'�9�K�]�o���X��  �Q_�S_\A�TBCKCTL.TM����ҟ����.�[INI�AeV~�SMESSAG!P�/�Q�@SQD�ODGE_D[P$VUb��O_�q��SPAUS�͠ !��K , 	��@�Eѯߧ,		ɯ�� '��#�]�G���k��� ����ۿſ�ͤ���?TSK  ��o<��PUPDTh�-��d~�~�XWZD�_ENB-��J��S�TA,��A~ŎAXI�S�@UNT 2��EQP� 	 �sR �߫kR"0`� Q�H�Ƹ�* ��/d�U�+�>�)�� v�� g��� 6_0X �� 5�!,����Pߊ�����METrK24�-S P���@h�
@K�k�@�*�7����?�I$@7|���>&I>.��=��f5RI�$<��>&+����SCRDCFoG 1�E�Q' �)UR�߆�������o�*Q %Ys�0�B�T�f�x��� ����������`,�����G�QGR���r���k��NA�P�K	�Th_ED�+�1V�� 
 ��%-��EDTA-Y�Z�M�1cC����R��*�BA�otV��)�u2~�[\���o�Q��/Yk/�w3 J/��/��s/�/%/7/�/[/w4?�/c? �/�??�?�/?�?'?w5�?R?/Ov?�O@vO�?�?eO�?w6�O O�OBO��OB_�O�O1_�Ow7z_�O�__ ��_oU_g_�_�_w!8Fo��o��oo@�o!o3o�oWow9�o_�o��;��o0�o�#wCR}�_ *�<��]�p���_���k � NO_DE�Lw�GE_UN�USEu�IGALLOW 1�	�   (*SYSTEM*���	$SERV_�GR��*���REG�3�$U���*�NU�MX�}�k�PMU|ր��LAY�����PMPAyL,���CYC1o��l�˝�����UL�SU��l�̒��5��L�?�BOXOR=I\�CUR_,�k��PMCNV���,�10����T4�DLI��%�G�	*�PROGRA2�?PG_MI���F��AL¥�����B�*�$FLU?I_RESUЗX�b����������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯�������H��k LAL_OUT� �T�WD_ABORѐ��j�O�ITR_RTN�  st��O�N�ONSTO� z�� b�CE_RIA3_I��z�������FCFG ��
��s}��_P}A9�GP 1����Q>�P�$b�!�C�p����z�-C�C ��(��+C8��@��H�� �CX��`��h��p���x}�����
�������	�su?���HE��O�NFI��Y�3G_mPr�1�� �� ă�}��������3KPAUSfI�1`�� �� �C`1oU� ������/5/@/Y/k/Q/�/Mo�NFO 1`��� � 	�-��/�p� ��	��@��>�"���vm�´��B��������/��CQ�Ch�@C3���ux��B���1�C��,B��Ã��I�䮵9l�fw�80��O�����sw�COLL�ECT_���&A���~7EN z��ܚ2W1NDE�3�7eヂ1234567890�7�~rD����?�6ss
 ���q)9O^OD�8O JO�OE�|O�O�O�O�O �O/_�O__w_B_T_ f_�_�_�_�_o�_�_ �_Ooo,o>o�oboto`�o�o�o�6B�2�;� �=�2IO  �9�1yxy�as؅�/wTR�2!}�� Jy
�o�~> �">}�z���9_MkORr#
� �Up�C(�n/X��! X�p�^�������ʋ1�T �q$?�,C?,,��UpK�TqJrJ��P[2&�?"�+�a�s�����
R���t7���u�y���5����s ���9PD�B/�(7��dcpmidbg�]�v &o�:��nD�pI����m�  ��nG�毱��ï��.�6����mg�x�C�Ůfg����-ſ�`ud1:���z~'�DEF 'y(�Is)��c�buf.txt�g��.%�_MC8�)7�!sd�ō�7�*������|��|�Cz  B3A�� Cظ�B���0CCI<g_}6�CC��-�E��D]qe�D�J0?����D�I�Df����-F��FR���F@��Cܤ��F@��F[��U|ɰ����,|P��t7AUpH Up�H �H ��t
���� ќ@ Da � D�  E	�� D�@ ��;��| Fp F"�� G=�fF���G'i�-G�>�Gg� G�K  H�<=H�&HyMc���  >�33 ' `C/��n)��F�5YT娂��A��|�=L��<#�� �Vq����ξ��RS�MOFST %x8ʝ/�&P_T1���DE -3�����q��Tq;�������?���<��;��EST2�+8�PR�2.a?����+C4���|��Up���������C��B�f��C����H��Up:d� ���T_~2�PROG ����%x�V$INU?SER  �5(�$KEY_TBL�  �"�	
��� !"#�$%&'()*+�,-./�7:;<=>?@ABC2��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������0�������������������������������������������������������������q* L�CKt��&t ST�AT���_AUT/O_DO�6���GIND�4�}1R����T27/�STqO@/� TRL, �LETE�7~*_�SCREEN �?�kcsc��2Uo MMENU� 1/.� < ED?[�/?J?ճ '?M?�?]?o?�?�?�? �?�?�?O:OO#OpO GOYO�O}O�O�O�O�O �O$_�O_Z_1_C_i_ �_y_�_�_�_�_o�_ �_oVo-o?o�ocouo �o�o�o�o
�o�o@ )vM_��� ����*���9� r�I�[������ޏ�� Ǐ�&����\�3�E� ��i�{���ڟ��ß��Ϲ�#_MANUAyLs/�!DBCO �RIG�'�/�_E7RRL2 0��a�aN�����ǯ P��NUMLI;�Z!�����
P�PXWO_RK 11�����'�9�K�]�o��DBwTB_�! 2���ç����DB__AWAYX�a�/GCP ��=E�ö�_AL;��òT�Y�r �%��I�_r� 1}3#� , 
�`T��B�ω�_M �I��Ѽ@����ON�TIM�'���ɼ���
�$�MO�TNEN��z$�R�ECORD 19Ξ� ��ψ�G�O�O�=߈�Ҳ{ߍ� �߱�Hع���O��s� (�:�L����߂��ߦ� ������� ���$��� H���l�~�������� 5���Y� 2D�� h��������� U
y�Rdv ����?�/ /*/�N/9/G/�/� �/�/�/;/�/�/q/&? �/J?\?n??}?�?? �?7?�?�?O�?�?FO �?jO�?�O�O�O�O_O �OWO_{O0_B_T_f_��OòTOLERE�NCдB��ްL���P�CSS_C�NSTCY 2:J����i_���_ �_�_oo'o9oKoao oo�o�o�o�o�o�o�o��o#�TDEVI�CE 2;�[ ��vu���������*��ϭSHNDGD <�[��Cz|{�TLS 2=]}<�����Џ�����>��RPA?RAM >0� ���|��}�SLAVE� ?]�I�_CF�G @J�*�d�MC:\�PL%04d.CSV)�b�cџ�RA ��CH�o�o�*��F��w�*�6�c�s�xa�`��JPѓ��|頪�r�_CR�C_OUT A�]}��.�_NOCO�D~�B0���SG�N C&��&j���20-A�PR-21 23�:42�*�0�9-FEB-18? 11:06��v LIX�v��r�*�s�Iu5��M��Þ��������VERSION -��V4.2.1�0��EFLOGI�C 1D�[ 	��+�ɘ�!���PROG_ENB��e�A�ULS�� �d��_ACCL{IM���������WRSTJNaT���*��MOJ������INIT cE�Z&�*� ��wOPTy� ?	�����
 	R5�75*�+�740�6J1�71�5�[�1U��21ԋ����TO�  ݉����V.��DEX��d��Hp���PATH ۦ��A\��9�K���[HCP_CLN�TID ?Ѷ��� ��"S��QI�AG_GRP 2�J�� Q� 	 @K��@G�?����?l��>��������Q �������P)��?�b�?�PT�i�^?�V�m?Sݘ���f403 6789012345{������� ��s���@nȴ@i��#@d�/@_��w@Z~�@U/�@O�@I��@D(���𷡋@���p����PAe�P�P�B4��jp��ط�
��1���-@)hs�@$��@ bN�@��@�����@�D@+����������	 ���R��@N�@I�@D��@>�y@9���@4� .v�@(��@"�\P�bt��L��@Gl�@BJ�@<z�@6��0��`@*� $N?�@���� $=q@����F@|��@33@��R@-?����?��`?�+hz����Y"�J�-@&��@N���!�?�?� � �//*/</�-�/ ?�/&?8?�/?Z?�? ^?�?�?@?R?�?�?O �?4OFO�?VO����@9�Q�i @��V���AY����?��z��A��5AF��A4��@��L4�R��A��@�p]� R�Q�R-P�P��@�� ��Ah���=H�9=Ƨ�=�^5=�>P��>���o=�,d_�,P�� ���C��<(;�U\� 4���ඨ_����A@��? ��pO�_xM�_o0o�� �T<ofo ovo�o~o�o��o|I>��y�b��R=���=���zq���G�G��� � ��!�!��NUt@�T��V���uB�� B��B��B%C�����~'����u���q�q6|䏁\�&���g���)PB�3pB�B A�@��"���m���<~��  5�-T��6�LT���o5���5����E���C�/�d�CO�ChA��l���r�ݏȏ���x�"�����C�3���u�lB���?H�� q�쏕�������ݟȟ� ���澺��Ƚ�ܷ�=��<��SxM��=���CT_CONFIG K�>m�eg7Ų��STBF_TTS��
YɈ�Ȱ��������MAU��N�N��MSW_CF\�L��  ��OCV7IEW��M�������A�S�e�w��� ����/�Ŀֿ���� ϭ�B�T�f�xϊϜ� +�����������,� ��P�b�t߆ߘߪ�9� ��������(��L� ^�p�����G��� �� ��$�6���Z�l�`~�������D�RC�	N(E��!P�����!�E4iX���S�BL_FAULT� O����GP�MSK���P�TD?IAG P`��q�o��o�U�D1: 6789?012345t�n���P*�Sew �������/ /+/=/O/a/s/2����R
B�/J�TR'ECP�
? )�+A>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^O�/�/�/�O��UMP_OPT�ION����ATR�袒��	�EPME����OY_TEMP�  È�3B��5P��TUN�I͠��5QܦYN_?BRK Q��?EDITOR�A�A�_�R_� ENT �1R��  ,�&ZAD15 �ADRA͠�_iH&STUDKW�_��_&-BCKE�DT-	o�^�R4 � %o7o�R3Oo�o�S2{o�o�S���o��M&STYL�E1�obo&PRgOG_�o<&}bs��P�t� ������/�A� (�e�L�������������ʏ܏� ��PMGDI_ST�Q�F5Q�}UNC;�1��� C�dO��v��N
�Nd�Oݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� �En���������ʑ�� ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@ߺ�g�q� �ߕߧ���������� �%�7�I�[�m��� ������������!� 3�E�_�i�{������� ��������/A Sew����� ��+=W�E s�������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?5?Oak?}?�?E? ��?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	__-_G?Y? c_u_�_�_�?�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7Q_[m� �_������!� 3�E�W�i�{������� ÏՏ�����/�I S�e�w��������џ �����+�=�O�a� s���������ͯ߯� ��'�A�3�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������9� K�U�g�yߋߥ����� ������	��-�?�Q� c�u��������� ������C�M�_�q� ���ߧ��������� %7I[m� ������! ;�EWi{���� ����////A/ S/e/w/�/�/�/�/�/ �/�/??3!?O?a? s?��?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O_ +?=?G_Y_k_!_�?�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	#_5_?Q cu�_����� ���)�;�M�_�q� ��������ˏݏ�� �-7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ����%�/�A� S�e��q�������ѿ �����+�=�O�a� sυϗϩϻ������� ���9�K�]�w��� �ߥ߷���������� #�5�G�Y�k�}��� �����������'�1� C�U�g��ߋ������� ������	-?Q cu������ �m��);M_y� �������/ /%/7/I/[/m//�/ �/�/�/�/�/�/!? 3?E?W?q{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O�O�O�O �O�O?�O+_=_O_i? __�_�_�_�_�_�_�_ oo'o9oKo]ooo�o �o�o�o�o�o�o__ #5G�os_}�� �������1� C�U�g�y��������� ӏ��o�-�?�Q� ku���������ϟ� ���)�;�M�_�q� ��������˯ݯ�	� �%�7�I�c�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ���������/�A� [�M�w߉ߛ߭߿��� ������+�=�O�a� s����������� ���'�9�S�e�o��� �������������� #5GYk}�� ������1 C]�gy���� ���	//-/?/Q/ c/u/�/�/�/�/�/I �??)?;?U_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�/�O_!_ 3_M?W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �O�o+E_;a s������� ��'�9�K�]�o����������ɏ�o �$�ENETMODE� 1TFu_�  �`�`��e�"��RRO�R_PROG �%��%�fe�r�@�TABLE  ���P��ß՟�@�SEV_NUM �  �	���@�_AUTO_?ENB  ,���=�_NO� U���!��  *U�]��]��]��]���+\�v�����6�F�LTR"�4�HIS���a�/�_ALMw 1V�� ��d]��`+��6�H� Z�l�~�����_��<�  ��[�"�պ��TCP_VER� !��!]���$�EXTLOG_R�EQ֦�-�'�SsIZ0�"�STKM��K��$�TOL�  �aDzޢ��A "�_BWD���������'���DI�� WFu�� ��a��STEP��������OP_D�Oo���FDR_G�RP 1X����d� 	пm�"�^�n�&���c?���$,M�T� ��$ ������^ӳ���^�B���IB�ĂB���BcGA?���A�R1����A�3B\��B���AIG��As� A��� ����:�%�^�I��m�����  @� ��As�Y>(������`
 E��q 	�����}+�������?�*�c���@�  ��@�33@%�������@����L�����^�F@ ������������L��FZ!D�`��D�� BT���@�����?� y M��6���u���5�Zf5�ES�����'�R��� ����`�X�����2�x�FEAT?URE YFu���&�LR �Handling�Tool ��b�English� Diction�ary�4D S�t� ard��A�nalog I/�O#,gle S�hift?uto� Softwar�e Update�dmatic B�ackup�	�g�round Ed�it� �Came�ra:F>Com�mon caliOb UI��n���Monitor��tr� Reli�abS�DHCP���
Data A�cquis�%)iagnos�7?+�ocument �Viewe"''u�al Check Safety�~�hanced�4�
�%s� Fr���xt. DIO ��fiu$�'end.� Err Lt"	=J�'s9r5�  ����
FCTN Me�nu� v##[7TPw InJ0facq5�GigE�>�5��p Mask Ekxc� g�'HT�0�Proxy Sv��$�6igh-Spe� Ski��6m ~� mmunic�7onsHurh0J0�:/;�2conne�ct 2:Hncr�0stru8Ja@�e�!� Jt%�KA�REL Cmd.� L�0ua�8�CR�un-Ti� Enyv�HK0el +��s�S/W�License�#�,0�Book(Sys�tem)�
MAC�ROs,�2/Of'fseZUH� w�8/"PMR �s.M�}M@!l�,Mec_hStop�1tQ@DY"Ui2V�Vx� �7�L^odTwiGtch�_aSh!.BV�[OptmoaS�0�fi�^aVg0GUulti-T�0��	PCM funkG:�ia�Ptiz~h�g�oV$RegiPr,@�fri� F�k�f�8Num Sel��U�i�  Adju�@�n qV1}tat�u�aI�*�RDM� Robots�cove�uea�v`� Freq AwnlyGRem�P��!n�u�rSer�vo� �P�SNPgX b�B[SN�0�Cli�!�WLi#br(��  �T:���vo�@th0ssag~e�� l5Q&��/I�=��MIL�IB����P Fi�rmu��Ph3Acyc��TPTX4/��eln5PǏ����1U��orquTi�mula!�E�u�PPa�A���!!c�&�0ev.��mr�i� �USR �EVNTğ֐ne�xcept� �pn��#ѕ�(@VC�rBB�XVU 6��G�4:�A�S�SC�y�gSGE����UI&?Web Pl`vǮ��q0O��0�$�!?6ZDT ApplD��
iP0a!�:� �Grid�qpla�y=����W�R-�.���h!N��B^P}2�00iV4+sciyi�1rLoad� �Upl���f@I�gPat�V�ycS`�B�`��� \6RL���� ۩�5MI Dev�@ (�qR�f�?��gsswo!�_�64MB DRA9MM���FRO�Ͼgell:�sh�D�#�c.k �rp��5�tySs
r7̬r'`.?+�p�!"=-o�� 2�a5por�t�.�p�r q�-T�1 �{]P��No� m�pc$筴OL��Sup��Fa�h?OPC-UA�l�#T �2eϓ�S0�0croa|�s:����~����uest�uS:��e2texV��u1p�1�#��PP�00�oVirt�!�sR��stdpnÛ�� �SWIMEST Mf F0������ �����������  MDVpz�� ����
I @Rlv���� ��///E/</N/ h/r/�/�/�/�/�/�/ ???A?8?J?d?n? �?�?�?�?�?�?O�? O=O4OFO`OjO�O�O �O�O�O�O_�O_9_ 0_B_\_f_�_�_�_�_ �_�_�_�_o5o,o>o Xobo�o�o�o�o�o�o �o�o1(:T^ ��������  �-�$�6�P�Z���~� ������Ə����)�  �2�L�V���z����� ������%��.� H�R��v��������� ����!��*�D�N� {�r����������޿ ���&�@�J�w�n� �ϭϤ϶�������� �"�<�F�s�j�|ߩ� �߲���������� 8�B�o�f�x���� ���������4�>� k�b�t����������� ��0:g^ p������	  ,6cZl� �����/�/ (/2/_/V/h/�/�/�/ �/�/�/?�/
?$?.? [?R?d?�?�?�?�?�? �?�?�?O O*OWONO `O�O�O�O�O�O�O�O �O__&_S_J_\_�_ �_�_�_�_�_�_�_�_ o"oOoFoXo�o|o�o �o�o�o�o�o�o KBT�x��� ������G�>� P�}�t���������� �����C�:�L�y� p����������ܟ� ��?�6�H�u�l�~� �������د��� ;�2�D�q�h�z����� ��ݿԿ� �
�7�.� @�m�d�vϣϚϬ��� �������3�*�<�i� `�rߟߖߨ������� ���/�&�8�e�\�n� �������������� +�"�4�a�X�j����� ������������' 0]Tf���� ����#,Y Pb������ ��//(/U/L/^/ �/�/�/�/�/�/�/�/ ??$?Q?H?Z?�?~? �?�?�?�?�?�?OO  OMODOVO�OzO�O�O �O�O�O�O_
__I_ @_R__v_�_�_�_�_ �_�_oooEo<oNo {oro�o�o�o�o�o�o A8Jwn �������� �=�4�F�s�j�|������̍  OH551���2�oR782�50��J614�ATU]P�545�6��VCAM�CUI�F�28H�NREv�52;�R63��SCH�DOCVCSU�869z�0�EIOCl��4��R69;�ES�ET$�:�J7:�R{68�MASK腯PRXYT�7�OCO�3$������m37�J6
�53���He�LCH�OP�LG$�0O�MHCuR �S��MATk��MCS#�0��55��MDSW�B�OPB�MPRC���s�]0�PCMS�5J�������s�51/�5u1{�0/�PRS697�FRDG�FwREQ�MCN�{93�SNBAx�^f�SHLB�M
�t����2�HTC#��TMIL􈳖TP�A˖TPTX<�EL۶����8�����wJ95_�TUTC�wUEV�UEC�wUFRG�VCC���OǦVIPG�CS�Ck�CSGk���I��WEB#�HTTf#�R6v���CG6�{IG�IPGS\��RCG�DGB�H7�5/�R7�Ry�Rk66O�2O�R6�WR55��4��5���D06�F�CL9I3�.�CMS˖0�n#�STY��TO7�q7��t�_�ORSǦt��M��NOM˖�OL�$���OPI^s�SEND�L��Sy�ETSsּ�SǻCPk�FVR˖I{PNG�Gene� È6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p�����	  ?H551���2�
R782�5�0�	J614�	AwTUP545�6�	VCAM�	C�UIF28lN�RE�
52[R6�3�SCH�	DO�CV�CSU�
8�690+EIOuC�4R69[�ESET<ZJ7�ZR68�
MAS�K�	PRXY|7.�
OCOL,3<�X 3�*J65u3�H�,LCH�*�OPLG<0�*M�HCR�*SJ;MA]T�MCS;0[+{55+MDSW�;v�+OP�+MPR�*t��,0PCM{�5KX +X0�+51�K51[L0KPR�SK+69�*FRD�kFREQ�
MC�N�
93SNByA��+SHLB�J�M[��<2HT=C;TMIL���TPA*TPTXF\ZEL�JX0�8
��
J95�TU�T�*UEVK*UE�C�*UFRkVCuC+lOk:VIPkZwCSC�ZCSG���I�	WEB;H�TT;R6��\C�G�kIG�kIPGmS�jRCkZDG�+�H75KR7:+R�YLR66�,2�*R]6�R55k|4�[]5�{D06+F�|�CLI�<JCMS�*�p;STY[kT�O�k7���OR�Sk:x M�LNO�M*OL�;�0�O{PI�jSEND�
uL:kSY�ETS�j� {[CP�FVR�*IPNkZGene��R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt������� ST�D�LANG ��	'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_�__q_�ZRBT�OPTN�_�_�_�_�_DPN�oo *o<oNo`oro�o�o�o��o�o�o�oted ��>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P bt������ �(:L^p ������� / /$/6/H/Z/l/~/�/ �/�/�/�/�/�/? ? 2?D?V?h?z?�?�?�? �?�?�?�?
OO.O@O ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8oJo\ono�o �o�o�o�o�o�o�o "4FXj|�� �������0�B�  �K�i�{��������Í99ʅ��$FEAT_AD�D ?	��������  	ǈ��,�>�P�b� t���������Ο��� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ �&�8�J�\�n����� ������������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O�O�O�O�O�DEM�O Y��   ǈ1]'_9_f_ ]_o_�_�_�_�_�_�_ �_�_,o#o5oboYoko �o�o�o�o�o�o�o�o (1^Ug�� ������$�� -�Z�Q�c�������Ə ��Ϗ�� ��)�V� M�_���������˟ ����%�R�I�[� ���������ǯ�� ��!�N�E�W���{� ������ÿݿ��� �J�A�Sπ�wω϶� �Ͽ��������F� =�O�|�s߅߲ߩ߻� �������B�9�K� x�o��������� ����>�5�G�t�k� }������������� :1Cpgy� ���� �	6 -?lcu��� ����/2/)/;/ h/_/q/�/�/�/�/�/ �/�/?.?%?7?d?[? m?�?�?�?�?�?�?�? �?*O!O3O`OWOiO�O �O�O�O�O�O�O�O&_ _/_\_S_e_�_�_�_ �_�_�_�_�_"oo+o XoOoao�o�o�o�o�o �o�o�o'TK ]������� ���#�P�G�Y��� }���������׏�� ��L�C�U���y��� ����ܟӟ��	�� H�?�Q�~�u������� دϯ����D�;� M�z�q�������Կ˿ ݿ
���@�7�I�v� m�ϙϣ�������� ���<�3�E�r�i�{� �ߟ����������� 8�/�A�n�e�w��� ����������4�+� =�j�a�s��������� ������0'9f ]o������ ��,#5bYk �������� (//1/^/U/g/�/�/ �/�/�/�/�/�/$?? -?Z?Q?c?}?�?�?�? �?�?�?�? OO)OVO MO_OyO�O�O�O�O�O �O�O__%_R_I_[_ u__�_�_�_�_�_�_ oo!oNoEoWoqo{o �o�o�o�o�o�o JASmw�� �������F� =�O�i�s�������֏ ͏ߏ���B�9�K� e�o�������ҟɟ۟ ����>�5�G�a�k� ������ίůׯ��� �:�1�C�]�g����� ��ʿ��ӿ ���	�6� -�?�Y�cϐχϙ��� ���������2�)�;� U�_ߌ߃ߕ��߹��� �����.�%�7�Q�[� ������������ ��*�!�3�M�W���{� ��������������& /IS�w�� �����"+ EO|s���� ���//'/A/K/ x/o/�/�/�/�/�/�/ �/??#?=?G?t?k? }?�?�?�?�?�?�?O OO9OCOpOgOyO�O �O�O�O�O�O_	__ 5_?_l_c_u_�_�_�_ �_�_�_ooo1o;o ho_oqo�o�o�o�o�o �o
-7d[ m������� ��)�3�`�W�i��� ����̏ÏՏ���� %�/�\�S�e������� ȟ��џ�����!�+� X�O�a�������į�� ͯ�����'�T�K� ]�����������ɿ�� ����#�P�G�Yφ� }Ϗϼϳ��������  �+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� �����	- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?m? ?�?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O__ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o������� ��#�5�G�Y�k�}� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-� ?�Q�c�u��������� ϯ����)�;�M� _�q���������˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߱����������� /�A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O��O_Y   XQ/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_
QPX3_E_W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������ ���/�A�S�e�w� ��������я���� �+�=�O�a�s����� ����͟ߟ���'� 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ����������	���$FEAT�_DEMOIN [ ԀK��!�}3�INDEX@��Oш3�ILEC�OMP Z�;����N�.��w�SETUP2 �[������  N ��t�_A�P2BCK 1\~��  �)�D����%���!��� �H����t���'� ����]�����(��� L���p������5��� ��k� ��$��1Z ��~��C�g ��2�Vh� ��?��u
/ �./@/�d/��/�/ )/�/M/�/�/�/?�/ <?�/I?r??�?%?�? �?[?�??O&O�?JO �?nO�OO�O3O�OWO �O�O�O"_�OF_X_�O |__�_�_A_�_e_�_ o�_0o�_To�_ao�o o�o=o�o�oso�o ,>�ob�o��' �K�o�������P�� 2��*�.VR�g��p*�j����s�����uQ�P�C��pFR6�:֏���;�ʋT _�_�q� �\���B�,�<���v*.FT��"�q	������C�қSTM c�l�w���d����piP�endant POanel��қH�������该�3�L�ӚGIFV�����l�)�;�пӚJPGڿϋ�`𿭿��T�ˊJS^�ć��p�u�2�%
�JavaScri3pt��޿CS�������ϵ� %Ca�scading �Style Sh�eets7ߩp
A�RGNAME.D)Tf��|��\z�8�К��Ի�g���DISP*�ߔߎ���>����0�?���	PANgEL15��%�� ���ﵯǯu�2���@�������o�z�3;�������L�^���z�4 ��%������wr��TPEINS.X3ML~�:\�P�bCustom Toolbar����PASSWOR�DC�~FRS:�\� %Pa�ssword ConfigW��4�/�ԝ[U�/q� �䘯���/�b_/v���/%J(�/g/y/?'2T/=?H(+? �/�/�?��?�/U5�?o?�?O'3\?EOH( 3O�?O�O���O�?]E �OwO�O_'4dOM_ H(;_�O_�_�_�O eU�__�_&o�Jo� no���o3o�oWo�o �o�o"�oFX�o| ��A�e�� �0��T��M���� ��=�ҏ�s����,� >�͏b�񏆟�'��� K���o�ٟ���:�ɟ ^�p�����#���ʯY� �}������H�ׯl� ��e���1�ƿU���� �� ϯ�D�V��z�	� ��-�?���c��χ��� .߽�R���v߈�߬� ;�����q���*�� ��`��߄��}��I� ��m�����8���\� n����!���E�W��� {���	F��j�� ��/�S��� �B��x��+��a�,�$�FILE_DGB�CK 1\������� < �)
SU�MMARY.DG�/�]MD::/z/��Diag S?ummary{/([CONSLOGp/�S/e!�/�/�!Co�nsole lo�g�/�\TPACC�N�/Y?%A?~?�%�TP Accou�ntin ?�Y@6�:IPKDMP.'ZIP�?�
�?O��%�0ExceptgionO�*�_�\O�bQJO�_1F�R DT Fil�es�O�<f MEMCHECKt?�/i/�_1Memor?y Data_��
l�)	FTAP�/f_�Oj_W1wmme`TBD�_��L >I)ETHERNET�_��A�_o�!Ethernet 0?figura&O�~}QDCSVRF�_pm__�oQ%]`� verify �all�o�M.=cXeDIFF�ovo��o P%�hd�iff�g�A]`CHG01�o���a5��b- `y2 ��&�1��gr�3����� �<�я`�VTRNDIAG.LS֏Ї���.�!Q� O�pe>c Log ~�!nostic����)VDEV�DA}O������aVisQ�D�eviceX�e�IMG��?����4�7�=ʔImag֟c�7UP{�ESz��?FRS:\z��O�@Updates� List����"�FLEXEVEANo�%�>��a� UIF Ev�Q�U�?�  ,�sz�)
PSRBWLOD.CMj���������0PS_RO�BOWEL�_�>*�HADOW4���+�D�SShad�ow Chang��O��a��RCMERR<�!�3����S��CFG �ErrorАta�ilk� �|�B��SGLIB��ЧϹ�N�!Q� S�t?`_�����):�ZDU_��7���nWZDT�adn�z���NOTIbo�߽�R�UNot�ific?b��t��{AGXbGIGE���/�A���]�GigExZ�d��N�A�� -��Q��^������ :�����p���); ��_����$�H �l��7�[ m�� ��V� z/!/�E/�i/� v/�/./�/R/�/�/�/ ?�/A?S?�/w??�? �?<?�?`?�?�?O+O �?OO�?sO�OO�O8O �O�OnO_�O'_9_�O ]_�O�__�_�_F_�_ j_�_o�_5o�_Yoko �_�oo�o�oTo�oxo �oC�og�o� �,�P���� �?�Q��u����(� ��Ϗ^�󏂏�)��� M�܏q������6�˟ ݟl����%���2�[� �������D�ٯh� �����3�¯W�i��� �����@����v�� ��/�A�пe����ϛ� *Ͽ�N����τ�ߨ� =���J�s�ߗ�&߻� ��\��߀��'��K� ��o����4���X� �����#���G�Y��� }������B���f��� ��1��U��b� �>��t	��$FILE_F�RSPRT  ���� ����$MDON�LY 1\8�  
 ��{� �������/ //�S/�w/�//�/ </�/�/r/?�/+?�/ 8?a?�/�??�?�?J? �?n?OO�?9O�?]O oO�?�O"O�OFO�O�O |O_�O5_G_�Ok_�O �_�_0_�_T_�_�_�_�o�_Co�_Poyo"VISBCKV@e*.VD�o�o8`�FR:\�`ION\DATA\�o�[b8`Visi�on VD file�oo>Pfot ^o�'��]�� �(��L��p��� ��5�ʏ܏�� ���$� ��5�Z��~������ C�؟g�������2��� V�h�#������?��� �u�
���.�@�ϯd��󯈿�)���LU�I_CONFIG7 ]8�aɻ� $ ��[{ 8 �2�D�V�h�zψ��|x���������� ��
ܠ�-�?�Q�c�u� ߆߽߫������ߊ� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi ����� �~/ASe ������h� //+/=/O/�s/�/ �/�/�/�/d/�/?? '?9?K?�/o?�?�?�? �?�?`?�?�?O#O5O GO�?kO}O�O�O�O�O \O�O�O__1_C_�O g_y_�_�_�_�_X_�_ �_	oo-o�_>ocouo �o�o�oBo�o�o�o )�oM_q�� �>�����%� �I�[�m������:� Ǐُ����!���E� W�i�{�����6�ß՟ �������A�S�e� w��� �����ѯ��� ���+�=�O�a�s��� �����Ϳ߿�Ϛ� '�9�K�]�oρ�ϥ� ���������ϖ�#�5� G�Y�k�}�ߡ߳��� �����ߎ��1�C�U�(g�y�	���x�����$FLUI_D�ATA ^���������RESULT� 2_���� ��T�/wi�zard/gui�ded/step�s/Expert ��"�4�F�X�j�|��������������C�ontinue �with G��ance��1CU gy������� ��-����0 ������6$���ps�o �������� /#/5/���\/n/�/ �/�/�/�/�/�/�/?�"?4?F>$(:Jrip�X�?�? �?�?OO*O<ONO`O rO�OC/�O�O�O�O�O __&_8_J_\_n_�_@�_Q?c?�_�?EJ��TimeUS/DST�_"o4oFoXo jo|o�o�o�o�o�o��?Enabl
 .@Rdv��P������ `�_��_�_f24o r���������̏ޏ�� ��&��o�o\�n��� ������ȟڟ���� "�4����)�;�M�zon
`7�ʯܯ�  ��$�6�H�Z�l�~����EST Ea��rn Stand������ӿ���	� �-�?�Q�c�uχ�� ��t�f�x�:|���acces�? �+�=�O�a�s߅ߗ�Щ߻�������ne�ct to Network���%� 7�I�[�m�����(����ȘB��Ϻ���ϊ�!��`Int�roduction��t����������� ����(�OL^ p������� $5�_�P�*����VEditor5����
//�./@/R/d/v/5 T�ouch Pan�el � (re�commen�P) �/�/�/�/�/?#?5? G?Y?k?}?�̬P�^��?��  �s/Reg`�O%O7OIO [OmOO�O�O�O�O6�EuropM�__ &_8_J_\_n_�_�_�_��_�_�_ B�z���?o�?�?��EU �_no�o�o�o�o�o�o �o�o"��C���B�an CeX�al ,ew�����@����+��V�L� o	oo-o?o������ Ώ�����(�:�L� ^�p�3������ʟܟ � ��$�6�H�Z�l� ~�:��QKY�k�}���>��/currNp�� �,�>�P�b�t�����𪿼�ο��14-F�EB-18 05?:03 PMԿ� �/�A�S�e�wωϛ��Ͽ���:�7�����pį֯���Yea� j�|ߎߠ߲�����������2018(�Q�c�u������������)� y
���  ���f�(�:���Month+����������,>Pbt��2 |������  2DVhz9�K���S\�n�������Day/$/6/H/Z/l/�~/�/�/�/�/��14�/�/	??-???Q? c?u?�?�?�?�?�?����O����HouY�fOxO�O�O�O��O�O�O�O__�5 $_J_\_n_�_�_�_�_ �_�_�_�_o"o�?�� Obo$O6O��inute'o�o�o�o�o );M_q�3x������ 
��.�@�R�d�v�5o��To��xo�o��AM����1�C�U�g� y����������)��� ��'�9�K�]�o����������ɯ��������Ϯ���ҏ�NetMethodϯ a�s���������Ϳ߿����0�Not� configureO�R�d�vψϚ� �Ͼ���������%�������!���� �߬߾��������� *�<�N�`�r� �ߗ� �����������'� 9�K�]�o�����b�L�Xߺ�|����� );M_q��� �x���%7 I[m���� ������/��3/E/W/ i/{/�/�/�/�/�/�/ �/?�?A?S?e?w? �?�?�?�?�?�?�?O O�:O�^O /�O�O �O�O�O�O�O__'_ 9_K_]_o_�O�_�_�_ �_�_�_�_o#o5oGo Yoko*O�oNO�orO�o �o�o1CUg y�����_�� 	��-�?�Q�c�u��� ������|oޏ�o��o Ə;�M�_�q������� ��˟ݟ����7� I�[�m��������ǯ ٯ����Ώ0��T� f�*�������ÿտ� ����/�A�S�e�$� �ϛϭϿ�������� �+�=�O�a� �j�D� �߸�z�������'� 9�K�]�o����� v��������#�5�G� Y�k�}�������r߼� ����
��1CUg y������� 	��-?Qcu� ������/�� ������\/�/�/�/ �/�/�/�/??%?7? I?[??�?�?�?�? �?�?�?O!O3OEOWO iO(/:/L/�Op/�O�O �O__/_A_S_e_w_ �_�_�_l?�_�_�_o o+o=oOoaoso�o�o �o�ozO�O�O �O' 9K]o���� �����_�5�G� Y�k�}�������ŏ׏ �����o.��oR� y���������ӟ��� 	��-�?�Q�c�t��� ������ϯ���� )�;�M�_����B��� f�˿ݿ���%�7� I�[�m�ϑϣϵ�t� �������!�3�E�W� i�{ߍߟ߱�p��ߔ� �߸���/�A�S�e�w� ������������ ��+�=�O�a�s����� ������������$ ��HZ����� ����#5G Y�}����� ��//1/C/U/ ^8�/�/n�/�/�/ 	??-???Q?c?u?�? �?�?j�?�?�?OO )O;OMO_OqO�O�O�O f/�/�/�O�O�/%_7_ I_[_m__�_�_�_�_ �_�_�_�?!o3oEoWo io{o�o�o�o�o�o�o �o�O�O�O�OP_w �������� �+�=�O�os����� ����͏ߏ���'� 9�K�]�.@��d ɟ۟����#�5�G� Y�k�}�����`�ůׯ �����1�C�U�g� y�������n������� ���-�?�Q�c�uχ� �ϫϽ������ϲ�� )�;�M�_�q߃ߕߧ� �����������"�� F��m������� �������!�3�E�W� h�{������������� ��/AS�t 6�Z���� +=Oas�� �h����//'/ 9/K/]/o/�/�/�/d �/��/��/#?5?G? Y?k?}?�?�?�?�?�? �?�?�O1OCOUOgO yO�O�O�O�O�O�O�O �/_�/<_N_Ou_�_ �_�_�_�_�_�_oo )o;oMoOqo�o�o�o �o�o�o�o%7 I_R_,_v�b_� ����!�3�E�W� i�{�����^oÏՏ� ����/�A�S�e�w� ����Z�~ȟ� �+�=�O�a�s����� ����ͯ߯񯰏�'� 9�K�]�o��������� ɿۿ����П�D� �k�}Ϗϡϳ����� ������1�C��g� yߋߝ߯��������� 	��-�?�Q��"�4� ��XϽ��������� )�;�M�_�q�����T� ��������%7 I[m��b�t� �����!3EW i{������ ���///A/S/e/w/ �/�/�/�/�/�/�/� ?�:?�a?s?�?�? �?�?�?�?�?OO'O 9OKO\?oO�O�O�O�O �O�O�O�O_#_5_G_ ?h_*?�_N?�_�_�_ �_�_oo1oCoUogo yo�o�o\O�o�o�o�o 	-?Qcu� �X_�|_��_�� )�;�M�_�q������� ��ˏݏo�%�7� I�[�m��������ǟ ٟ럪��0�B�� i�{�������ïկ� ����/�A� �e�w� ��������ѿ���� �+�=���F� �jϔ� V�����������'� 9�K�]�o߁ߓ�R��� ���������#�5�G� Y�k�}��NϘ�rϼ� �����1�C�U�g� y��������������� 	-?Qcu� ���������� ��8��_q��� ����//%/7/ ��[/m//�/�/�/�/ �/�/�/?!?3?E? (�?L�?�?�?�? �?OO/OAOSOeOwO �OH/�O�O�O�O�O_ _+_=_O_a_s_�_�_ V?h?z?�_�?oo'o 9oKo]ooo�o�o�o�o �o�o�O�o#5G Yk}����� ��_
��_.��_U�g� y���������ӏ��� 	��-�?�P�c�u��� ������ϟ���� )�;��\����B��� ��˯ݯ���%�7� I�[�m����P���ǿ ٿ����!�3�E�W� i�{ύ�L���p��ϔ� ����/�A�S�e�w� �ߛ߭߿����ߢ�� �+�=�O�a�s��� �������� ���$� 6���]�o��������� ��������#5�� Yk}����� ��1��:�� ^�J������ 	//-/?/Q/c/u/�/ F�/�/�/�/�/?? )?;?M?_?q?�?B� f�?�?�OO%O7O IO[OmOO�O�O�O�O �O�/�O_!_3_E_W_ i_{_�_�_�_�_�_�? �?�?�?,o�?Soeowo �o�o�o�o�o�o�o +�OOas�� �������'� 9��_
oo~�@o���� ɏۏ����#�5�G� Y�k�}�<����şן �����1�C�U�g� y���J�\�n�Я���� 	��-�?�Q�c�u��� ������Ͽ����� )�;�M�_�qσϕϧ� �����Ϝ�����"�� I�[�m�ߑߣߵ��� �������!�3�D�W� i�{���������� ����/���P��t� 6ߛ����������� +=Oas�D� �����' 9K]o�@��d� �����/#/5/G/ Y/k/}/�/�/�/�/�/ ��/??1?C?U?g? y?�?�?�?�?�?��? �O*O�/QOcOuO�O �O�O�O�O�O�O__ )_�/M___q_�_�_�_ �_�_�_�_oo%o�? .OORo|o>O�o�o�o �o�o�o!3EW i{:_����� ���/�A�S�e�w� 6o�oZo��Ώ�o��� �+�=�O�a�s����� ����͟����'� 9�K�]�o��������� ɯ�������� ��G� Y�k�}�������ſ׿ �����ޟC�U�g� yϋϝϯ��������� 	��-�����r�4� �߽߫��������� )�;�M�_�q�0ϕ�� ����������%�7� I�[�m��>�P�b��� ������!3EW i{������� �/ASew ���������� /��=/O/a/s/�/�/ �/�/�/�/�/??'? 8/K?]?o?�?�?�?�? �?�?�?�?O#O�DO /hO*/�O�O�O�O�O �O�O__1_C_U_g_ y_8?�_�_�_�_�_�_ 	oo-o?oQocouo4O �oXO�o|O~o�o );M_q��� ���_���%�7� I�[�m��������Ǐ �o菪o���E�W� i�{�������ß՟� �����A�S�e�w� ��������ѯ���� �؏"���F�p�2��� ����Ϳ߿���'� 9�K�]�o�.��ϥϷ� ���������#�5�G� Y�k�*�t�N����߄� ������1�C�U�g� y����������� 	��-�?�Q�c�u��� ������|ߎߠ߲� ��;M_q��� ������7 I[m���� ���/!/���� f/(�/�/�/�/�/�/ �/??/?A?S?e?$ �?�?�?�?�?�?�?O O+O=OOOaOsO2/D/ V/�Oz/�O�O__'_ 9_K_]_o_�_�_�_�_ v?�_�_�_o#o5oGo Yoko}o�o�o�o�o�O �o�O
�O1CUg y������� 	��,?�Q�c�u��� ������Ϗ���� �o8��o\������� ��˟ݟ���%�7� I�[�m�,�������ǯ ٯ����!�3�E�W� i�(���L���p�r�� ����/�A�S�e�w� �ϛϭϿ�~������ �+�=�O�a�s߅ߗ� �߻�z��ߞ� ���� 9�K�]�o����� �����������5�G� Y�k�}����������� ���������:d &������� 	-?Qc"�� ������// )/;/M/_/hB�/ �/x�/�/??%?7? I?[?m??�?�?�?t �?�?�?O!O3OEOWO iO{O�O�O�Op/�/�/ �/_�//_A_S_e_w_ �_�_�_�_�_�_�_o �?+o=oOoaoso�o�o �o�o�o�o�o�O �O�OZ_���� �����#�5�G� Y�o}�������ŏ׏ �����1�C�U�g� &8J��nӟ��� 	��-�?�Q�c�u��� ����j������� )�;�M�_�q������� ��x�ڿ������%�7� I�[�m�ϑϣϵ��� ������� �3�E�W� i�{ߍߟ߱������� ���ʿ,��P��w� ������������ �+�=�O�a� ߅��� ����������' 9K]�~@�d� f���#5G Yk}���r�� ��//1/C/U/g/ y/�/�/�/n�/��/ ?�-???Q?c?u?�? �?�?�?�?�?�?O� )O;OMO_OqO�O�O�O �O�O�O�O_�/
?�/ ._X_?_�_�_�_�_ �_�_�_o!o3oEoWo O{o�o�o�o�o�o�o �o/AS_\_ 6_��l_���� �+�=�O�a�s����� ��ho͏ߏ���'� 9�K�]�o�������d v�����#�5�G� Y�k�}�������ůׯ ������1�C�U�g� y���������ӿ��� 	�ȟڟ�N��uχ� �ϫϽ��������� )�;�M��q߃ߕߧ� ����������%�7� I�[��,�>Ϡ�b��� �������!�3�E�W� i�{�����^߰����� ��/ASew ���l������� +=Oas�� �����/'/ 9/K/]/o/�/�/�/�/ �/�/�/�/� ?�D? k?}?�?�?�?�?�? �?�?OO1OCOUO/ yO�O�O�O�O�O�O�O 	__-_?_Q_?r_4? �_X?Z_�_�_�_oo )o;oMo_oqo�o�o�o fO�o�o�o%7 I[m��b_� �_���o!�3�E�W� i�{�������ÏՏ� ���o�/�A�S�e�w� ��������џ���� ��"�L��s����� ����ͯ߯���'� 9�K�
�o��������� ɿۿ����#�5�G� �P�*�tϞ�`����� ������1�C�U�g� yߋߝ�\��������� 	��-�?�Q�c�u�� ��X�j�|ώ����� )�;�M�_�q������� ����������%7 I[m���� ���������B� i{������ �////A/ e/w/ �/�/�/�/�/�/�/? ?+?=?O? 2�? V�?�?�?�?OO'O 9OKO]OoO�O�OR/�O �O�O�O�O_#_5_G_ Y_k_}_�_�_`?�_�? �_�?oo1oCoUogo yo�o�o�o�o�o�o�o o-?Qcu� �������_� �_8��__�q������� ��ˏݏ���%�7� I�m��������ǟ ٟ����!�3�E�� f�(���L�N�ïկ� ����/�A�S�e�w� ����Z���ѿ���� �+�=�O�a�sυϗ� V���z����ϲ��'� 9�K�]�o߁ߓߥ߷� �����߬��#�5�G� Y�k�}�������� ��������@��g� y��������������� 	-?��cu� ������ );��D��h�T� ����//%/7/ I/[/m//�/P�/�/ �/�/�/?!?3?E?W? i?{?�?L^p��? �OO/OAOSOeOwO �O�O�O�O�O�O�/_ _+_=_O_a_s_�_�_ �_�_�_�_�_�?�?�? 6o�?]ooo�o�o�o�o �o�o�o�o#5�O Yk}����� ����1�C�oo &o��Jo����ӏ��� 	��-�?�Q�c�u��� F����ϟ���� )�;�M�_�q�����T� ��x�گ����%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ���ʯ,��S�e�w� �ߛ߭߿�������� �+�=���a�s��� �����������'� 9���Z��~�@�B��� ��������#5G Yk}�N��� ��1CUg y�J��n���� 	//-/?/Q/c/u/�/ �/�/�/�/�/�?? )?;?M?_?q?�?�?�? �?�?�?���
O4O �[OmOO�O�O�O�O �O�O�O_!_3_�/W_ i_{_�_�_�_�_�_�_ �_oo/o�?8OO\o �oHO�o�o�o�o�o +=Oas�D_ �������'� 9�K�]�o���@oRodo�vo؏�c�$FMR�2_GRP 1`���� ��C4  B�.�p	 �p�0���F@ F�E���Q�F���C��L��FZ!D�`��D�� BT���@���^�?� � �����6��������5�Zf�5�ESΑ^�A�3  ���BH��\�~�@�33@��	 ����@�Q���@�g�]�Q����<��z�<�ڔ=�7�<�
;;�*�<��^��8ۧ�9k'V�8��8����7ג	8(�� ~�����=�(�a�L�����w�_CFG a�T0���ӿ�|����NO �/
F0+� 0����RM_CHKTYP  �p	������ROMF�_MsINL��s��x�u�7�X�SSB���b�� ��Ϛu�����ϝ��TP_DEF_O/W  �t	��ǟIRCOMK�����$GENOVRD�_DOm��q*�T[HRm� dG�d0�o_ENB� 0ЯRAVC��c���� �>�����v����^����.� ���OU��i��3�.��.�< u�����,�z����sC�  D����l�d�$�@��B�/���1�m��ϑ�SMT���j��������$�HOSTC��1k������� kMC�t�����v  27.0z 1��  e�� BTfx�
0�������	anonymous 4FXj|�r���������)
/ /./@/R/�v/�/�/ �/�i/�/??*? <?N?����?�/�? ��?�?OO�/�?JO \OnO�O�?�O�/�O�O �O�O_S?�Ow?�?j_ �O�?�_�_�_�_�_+O oo0oBoTow_�O�O �o�o�o�o�o'_9_K_ ]__o5�_t��� ��_����(�K }o�op����������o 13�$�gH�Z� l�~������Ɵ؟� ���Q��D�V�h�z� ��Ϗ�󏥯���;� �.�@�R�d������� ������%���*� <�N�`ϣ���ǯ��ۿ �������&�i�J� \�n߀ߒߵ�7�����������"�o���EN�T 1l��� � P!��s�  v�a�������� ��
������?�d�'� ��K���o��������� ��*��Nr5� Yk����� 8�1n]�U� y����/4/� X//|/?/�/c/�/�/��/�/�/?�/B?:?QUICC0O?+?=?�?a41�?{?�?�?�a42�?�?�?>O!?ROUTER?OO�-O�O!PCJO�G�OjO!19�2.168.0.�10h?]3CAMP�RT�O�O!�E1�@_�FRTXO
__�}_C�NAME �!P�!ROBO��O�_S_CFG �1kP� ��Auto-s�tarted��FTP��a�Ϧ� Ao��eowo�o�o�oF� �o�o�o*o�oO as���r��_o o�'Io�<�N�`� r�5������̏ޏ� ���&�8�J�\�n�g� yϋϝ�鏿����� "�4�F�	�j�|����� ��՟W������0� B�������������� ҿ�����ݯ>�P� b�tφϩ�+ϼ����� ����Y�k�}�/ߑ� ��ſ�߸������߱� �$�6�H�k�l��ߐ� ���������-�?�Q� 2�e�V���z������� s�������
?��� ;dv������ �%�9[�<N` r�G����� �&/8/J/\/n/�/ ������//? "?4?F?X?/|?�?�? �?�?�/i?�?OO0O�BOTO�Z_ERR �m�Z\OlFPDU�SIZ  �0^�0��D>�EWR�D ?�U�!� � guest�6�O�O __$_�6_�TSCD_GR�OUP 3n�\ u�Q�9IFT|^w$PA|^OMP|^w |^_SH|^�ED�_ $C|^C�OMn@TTP_A�UTH 1o{K� <!iPen�danBWMn�[�2��q!KAREL�:*MoVohmKC�}o�o�ou`VISION SETfP�o�o�v!,rc P>hb�������~dCTRL Kp{M6��1
F��FFF9E3���$FRS:D�EFAULT[��FANUC W�eb Server[�I��"d�O�D��я�����+�jDW�R_CONFIGw qkU�B�c[�lAIDL_C_PU_PCz��1sB�� �� BH���MIN��sQ��GNR_IOuA�B�0�H���NPT_SIM�_DOӖݛSTAL_SCRNӖ� �ޚTPMOD�NTOL�ݛ��R�TY������` `E�NB�sS��OL_NK 1r{KxP ����ɯۯ������_MASTEҐy��5���SLAVE �s{KH D��S�RAMCACHE�/�A�"aO_CFGq�����UO�`����?CMT_OPz�ՒJǳYCLp���t�_ASG 1t`��A
 �6�H�Z� l�~ϐϢϴ����������� ��	�NUMj�CI
��IPn����RTRY_CN8ҿ���_UP_��A�����E ������]u)�  06������RCA_ACC� 2vk[  R��� 1q� � j� 6�� W6��0+�4�?4�� 9"��� �2D���BUF�001 2wk[=� �u��u0����u0�pi�u0_�n�)��8��UI��X��i��x��U��䘞䩞丞�Uɞ�؞������C	��� ����U�����������������������u0��Zx��U��!��0��A��UP��a��p���}����;@  ��Ӗ� ����������$��3��D���S��d��s����䓖�u0��l����Ɩ����s�2������ޤ�u ��t(������ ����������t� ����� ����� ��$�)��)�<�) �L�)�\�)�l�8)�|�K *����phȜ��� �������� ������������������" t� �� �  �% �- �5 �=  �E �M �U �]  "e �m �u �s�3���.��.�-� �@���.����.��� �.����.���.� �.��#�R%�3 �R�$<�K�R�$T�c �R�$l�{�R}��P� �P���P������ ���������� ���������R�� #i�#i�+#i� -;#i�=K#i�M[# i�] i�es#i�u����я�2xk[ 4�6�A��Q�P<�Pp�D�AՒ��HIS}��zk[ �� �2021-04-;21�V ��A �I/_A_S_e_w_�_�_x�_�_�XR��yX 	CT�_
oo.o@oRo`dovo�o�o���y��;  L[T�Q�18-02-27��_�o�o�o  T�c,>Pbt�{/LY�3�h5�o�@�������U�p*G�Y��sN�2�g1�A�������\��C����BXQ�``΄h�ބiC�D���΄��2��(�:�LM��@u�2���q����H<&q���F�:�p΄x@ބF��A�Q�A�΄5�΄�΄�����rL��u��`�M�_� q��FՂƐ݂�@��@�ђ�`ْ�@��������M� �O_Z: �M�_�q����� ����˿ݿ��_;�%� 7�I�[�m�ϑϣϵ�
�n;�@c�o����%�7�%p5  Z 8�c�u߇ߙ߇��� ������)�;�)�M� j�|�j�|�������ĉB�AdՀ��݀6�d������������ -
�@L�6Z�O�=�O� ����������Ɛ� ѐ�ⵠ������ P��ՠ�����	��� ���&�8�n���� ��݀��
���ѐ� ��*	�9�L� �&�Z�|�� �����/��� /T/f/x/�/�/�/�/�/�/�d����:/'?9?K?9���#v?�?�? �?�?�߾�?OO*O<ONO`O)�iO�O�O ����O�O�OŊ���@ ݂���@��@��~O
� BR�B_s_�Os��O�_ �_���_��4Xђ�P�� �P��
��P͢�Pբ�P ��P	��P�_oM�_ �o�o�o��$_o$o6o�Ho�;�I_CF�G 2{: H�
Cycle �Time�aB�usyDwIdylzr�tmin={=�qUpvv|q�Read�w�Dow�x�aR}qsCount|q�	Num qr�s��={��`�!�PR�OGWr|:D�0�u����������Ϗ�y%SDT_ISOLC  :�� �@~J23�_DSP_ENB�  �>#�IN�C }��e�A�   ?��=�̟�<#�
�j�:�o u������aX��ȟ�OBK�C,���uU��G_GR�OUP 1~�}< � �Pj�Cy.�П?Dxd�m��`Q������̯�� ���&�Dw��ڙ�G_IN_AUT�O�Q�#�POSR�E���KANJI�_MASK��t�K�ARELMON #:(��by�π�(�:�L�@~²O��V�X��nŉ����CL_Ld�NUM�0�����EYLO�GGING��?����U�F�LANGU�AGE :�
��DEFA�ULT �(LGfXq�V��r��d?�  8�pPu��`'6'  ��`�ۏ�;��
���(UT1:\\Ϧ� �ߵ����� �����!�8�E�W���(��#LN_D?ISP �M��x�������OCTOL���aDz@��f���GBOOK ��)�=z�qz�z�=  �ey�k�}���������`��5Ӱs����	-��t�*��/ُ`�+�_BUFF 2��O A�ev ꂒ�w���� �#,YPb� �������/���ZDCS � V�Y�n���#Dx^u�/�/�/�/6$IO 2�B+ cp�/cp@���/??*?>?N? `?r?�?�?�?�?�?�? �?OO&O8OJO^OnO��O�O�O�%ER_ITM��dD��O_#_ 5_G_Y_k_}_�_�_�_ �_�_�_�_oo1oCopUogo	��BSEV������FTYP����O�o�o�ovm��RS�T��4%SCRN__FL 2��-@��g/gy������TP�����b>�NGNAM,�`��
�2$UPS��GI�p��U�B�_L�OAD�G %� �%ZAD15��O�MAXUALcRM�¢� �U�9
��H�_PRM���� !���C����7������P �2�7� �V�	 �ol�W���{���Ɵ�� �՟���D�/�h� S�������¯���ɯ ۯ��@�+�d�v�Y� ������������߿� �<�N�1�r�]ϖ�y� ���Ϸ������&�	� J�5�n�Q�cߤߏ��� ��������"��F�)� ;�|�g�������� �������T�?�x� c����������������DBGDEF ��[!��_LDXDISA-��{�#MEMO_AP'��E ? �
 $x(�����������FRQ_�CFG ��6(A x'@�E��<[$d%m$�:������*�/� **:�����_x& ��+/"/4/a/X/j/ �/����/�@�/�/�/�/�',(�/>?�$,? i?P?�?t?�?�?�?�? �?OOOAO(OeOwO�^O�O��ISC 1� �� ����O�� )�O��2__V_�O�B�_MSTR ���myUSCD 1�o�N_�_J_�_�_o �_4oo1ojoUo�oyo �o�o�o�o�o�o0 T?xc��� ������>�)� N�t�_����������� ˏ���:�%�^�I� ��m�������ܟǟ � �$��H�3�l�W�i� ����Ư���կ��� �D�/�h�S���w���؛�Կj_MK'���]Y�$MLTA[RM&�-� 3" P�X� �METPUK Ȳ����YNDSP_ADCOLr�& }�oCMNT�� ���FN���τ�FST�LI���ǁP ���^'�G�Y?�IԆ�P�OSCF����PgRPM��Y�ST���1��[ 4Q#�
��ϱ�����׿� ������7��+�m�O� a��������������E�/��SIN�G_CHK  ���$MODA%��K���DEV� 	N
	MC}:��HSIZEK�Ȱ��TASK �%N
%$123456789  �2}�TRIG 1��[ l^`9n�=YP���5��~�EM_I�NF 1���`)AT&FVg0E0�+)�E0V1&A3&�B1&D2&S0�&C1S0=)�ATZ+fH@��:��bA�@/�'//K/]/  �/5GYk�/� ? 7/$?6?�Z??~?�? w?�?g/y/�?�/�/�/ 2O=?�/hO�?�OGOQ? �O}O�O�O
__�?@_ �?OO)O�_MO�_�O �_�_�Oo�_<oNo5o ro%_7_�o[_m__�o �_&]oJo� ;�����o��o �o�o�oX�|���� ��e֏�����0����NITOR�G� ?��   	?EXEC1˳s�U2y�3y�4y�5y�TC {�7y�8y�9˳t��rޔx�ޔ��ޔ ��ޔ��ޔ��ޔ��ޔ@��ޔ̒ޔؒޓ2�U2�2��2	�2�U2!�2-�29�2E�U2Q�3�3�3����R_GRP_S�V 1�  (�7���;=�/�";���������ɿN?�����
_Dς��9��ION_DB��|��ȱ  �q�fh�G��~� Ȱ����ΰ.ΰ/���&�N   1�ڿ����J��-ud1����υ��PL_NAME �!<��!�Default �Personal�ity (fro�m FD)����R�R2�� 1�L?6�LA�<��� d:҉ϛϭ� ����������+�=� O�a�s߅ߗߩ߻���������2��.�@� R�d�v���������<�����0�B� T�f�x����������$޲�����
���PJ\n�� ������" 4FX'9��� ����//0/B/ T/f/x/�/�/k}�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�>� H�6 H?�b H\����  �O1M�d C@PObMFO�O�G@ �=�|C�O�M�O�O C �H__ _2_ P_V_t_�_�f��_�\��E	`_�_o| o�Q:�oA`��@oRodovn A�  �i�O�o�Lޱ �o�k�O�o'9$�]H� �R�� 1�4ɴ��R@ �� &�<��p �@D�  �q?���s�q?��q�A�?�6Ez  �q����;�	l�r	 ��@�? 0ݰް�!� ��p� � �� �F��J���K ��J�˷�J� �J�4�JR�<g|�v�f0O���@�S��@�;fA6�A��A1�UA��X{�����=�N��f������T;f��X��ڀ���*  ��  ?�5��>��p��H��?��?����#�����ԏur`�f��q`{��g������i��V���(  �����Ȗt����	'� � ��I� � � ��e��:����(�È=����@����� <�!�� � �  ��qz���r�o�o��<��ү  '覵���@!�p@�a��@��@��@��-C�C"��"���B�pC%�����@�r�������n�������m;a;n�`@����D�u՟ҿ �������Q�c�E��Uŕ�� :�W � x�x?�ff0�O�Ϙ�*� �P����ˍ�8�����>����x��q����0�P�:�U�7�0�0���>��|���<2�!�<"7�<L���<`N<D��<��,h��ߴ��s���s ҈`?ff�f?��?&�аT@�T���?�`�?Uȩ?X� ᒩL����t,��t8� �wW�����ό�w�� ����������.��R���!�F�A��� =���)���M����HmN H[���G� F�� HZE~i��� ���� �oAK ��������)� ��/��%/7/�j/ U/�/y/�/�/��M��"�i��C�/?�/5? =8��??F??j?���ç�s��-M�BH�"��.��?,�[2�xY0X1�1@Iܔ=�@n�@���@: @l���?٧]�? ���%�n��߱���=�=�D��0OB@���@�oA�&{�C/� @�U�XO�+J8��
�H��>��=3�H��_�O �F�6�G���E�A5F�Į�E��O�@���fG��E���+E��EX���O�@>\�G��ZE�M�F�lD�
�p�O�? E_0_i_T_�_x_�_�_ �_�_�_o�_/ooSo >owobo�o�o�o�o�o �o�o=(:s ^������� � �9�$�]�H���l� ������ۏƏ���#� �G�2�W�}�h����� ş���ԟ���
�C� .�g�R���v������� �Я	���-��Q�<��u�`�r���fB(hA4g���h������3�ϩп��!�4 �{����!��0+#(�:��j�bT�f�1E���|�Ђˀ��Ϯ���P�����iP��P:�IVc߶�oߙ߄��ߨف����������9�$��"$<�N�� r�����v�H���&��e,�6�l�Z�|�����n)���������8F
  2� H�6�&H�,{�g\��&B�!�!�� B��0�0A� @ �/��$�3���l^pUgy����$0� �� ��� T�%
 ��//+/=/ O/a/s/�/�/�/�/�/��/^J� ��$�����4�$MR_�CABLE 2�>$� � V�UTP��@{ ?�0�F1�?0��0z B�z C[0{OM�`oB���{�0�#DG�l{??Q65  B�� T�O
�vr0���w5Ų~6q<�|�h�?�8� �� C� ]9h4��r0��2w��E~6�'N�?��?�*\0�� [@C�W@j27�(��{<��2I�/T3 �OR˰O�O�O�O�O_ �O�O"__*_�_�_`_ �_�_�_�_�_oA{+��_Qocouol�?op�o�o�ol�*�o�** 3OM }�%9��z{�0�3%% 23�45678901%7u "RFq{ [@� �{ {
�Lw�nnot s�ent �jzsW�,�TESTFECSALGRI��gkʝd�t��q
,�tG �P�{�"���'�9�K� 9�UD1:\mai�ntenance�s.xm�7��l����DEFA�ULT2GRP� 2�	z  p�$�  �%1�st mecha�nical chgeckL}{�6�#�>�G�H�$�r���������{�c�ontrolleAr��7��Ic��8�J�\�n���ϑMX���{"8��{ ȡϯH'�����*�<���Cٟn����������ҿ�����ϒC�ge�. battery���W�H	���ϖϨ������ϑSupp�ly greasXK���{��
�<A��g�s�H�Z�l�~����ϑ �cabl��߾�g�
7��� 0�B�T��ؑ+�����Q������������{ $��@�hoo�  �����������+�  O�a�s�)Zl~� ����'9  2DV���{ ����
//k@/ R/�v/��/�/�/�/ �/1/?U/g/<?�/`? r?�?�?�?�/�??-? OQ?&O8OJO\OnO�? �O�?�?�OO�O�O_ "_4_�OX_�O�O�_�O �_�_�_�_�_I_om_ _To�_xo�o�o�o�o o�o3oEoWo>P bt��o��o ���(�:���p� �_����ʏ܏� � O�$�6���Z���~��� ����Ɵ��9�K� � o�D�V�h�z���۟�� ����5�
��.�@� R���v�ůׯ����п �����g�<ϋ��� r����ϨϺ�����-� �Q�c�8߇�\�n߀� �ߤ������)�;��� "�4�F�X�j�ߎ��� �����������m� ��T���C�������� ����3�i�>�� bt������ /S(:L^p��	 T~�� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�?�OO0OBOTOfOxO � �?�  @� ��O�O��O��O__(_�;*H_** �� �@zO|_�_�_b_�_�_�_�_��!__ �_Ko]ooo1o�o�o�o oo%o�o#5o Ak}��o�oQ� ��E�1�C�U�� ��a�����ӏ�����	��e�w��
�$M�R_HIST 2���v�� 
 �\�$ 2345?678901����P�BR��9���� �����?�Q�c��,� ������t���ԯ�� ί;��_�q�(���L� ��˿��￦��%�ܿ I� �m��6ϣ�Z�����ϐ���[�SKCF�MAP  ��y��B������ONREL  ��v�.�6���EXCFENB�`�
,��y�FNC���r�JOGOVL�IM`�dv����K�EY`�����_�PAN_������R�UN����SFSPDTYP��k���SIGN`�r�T1�MOT��o��_�CE_GRP 1��.�~���O ��÷���a������ C�U��y�0�����f� ������	��-?& c����t� ���Mq�(�QZ_EDI�T]�(�Q�TCOM_CFG 1�$�a����� 
�__ARC_}�`����T_MN_MO�DE]���UA�P_CPL/��N�OCHECK ?�$� ��  �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�?�I�NO_WAITc_L\���NT���$�3���1_7ERR��2�$�6���OEOWOiO�L<юO��O�53 OC�#M|� 1q�f?"���A,:?x���k��µ�_B��z��<�� ?���_�O?�|7NBPARAMB�$���Fg�_pyW8ѫ_�[ = �� �_�_�S�_o(oo4o�^opoLo�o�o�kxW���o�l}_n#UM_RSPACE!���b�GQt�$OD�RDSP#_��O�FFSET_CAqR�_/�vDIS��sS_A3 ARK�]�OPEN_FILE�p_���cq�PTION_IO������M_PRGw %3z%$*A�lS��sWO�p����C쀄���ꂗ  ;�?֞��g��	 ��Ȟ�����4�dpRG_DSBL  n��.�J��sRIE�NTTO_���Cٴ>�-�A �rUT�_SIM_D��+ҋBdpVhpLCT ��=���O}��=d\�_PEX; �n��RAT;' d������pUP �m��pw���� �|>�L��$PAL�2���>`�_POS_CCH�p��`�ZP2����L6�LA�W����oѯ �����+�=�O�a� s���������Ϳ߿� ��'�9ϳ�2��h� zόϞϰ��������� 
��CW�4�F�X�j�|� �ߠ߲���������* AAs'�}I5�4�Z�BPG��������� ����&�8�J�\�n� ����a�s��������� "4FXj|� �������� 0BTfx��� ����///_�xW�Y/k-���c�� �/�+�/�/�'>->-�o?�/3?�'tP(7R? H?Z?l?�?�?�?�?&0`w��?L�D(4	`<?�6OHOZOA:�o�<�xO�O�O�O'0A�  �I!?�O�__ �]?>_)_b_M___�_��_�_u����O�1�������� ��$B@ ��؄��P @D��  a?�c�Q?�=�a=�D�  E�z0c�:�;�	l�&b	 �@�� 0�PP_` �
`�� � � ���b�PH0#H���G�9G��ģG�	{Gkf���GΈK/�o�l�P�C�1��`[�D	� D@ D7g��n�d���  ß5��>(p`�p4�(: B4��Bp{�!�=���O��R ��r'a�sW�Ao�R�ҧpߐ�p(�  ��p�����_$��U	'� �� B�I� ?�  ��E�F�=���f�x��߶� <_`�� � � ��ف��8�" b__�WN=���  'N�(��aOpC��`��`[pB`C�c5�G� ���@��i���~�m����G�MuAuN�@@=��*b 7e����4��X�C����������=�� :��a�tx?��ff�/į֯h� @��O�8=�3�A�>�׶q"a�J�pn�Px���uancnd؃�>������u<2��!<"7�<L���<`N<D?��<��,�o㿌�c� c^��@?offf?�?& ��K�@T�2�?��`?Uȩ?X�B�:銒�'d�I ev�g���Zd���� ���������6�!�Z� l�Wߐߢ�y��߱����aσυ���D���Hm�N H[��2G�� F��M��� �����������(� �%�^� _���K�� ���+���g�*< N�cu������Β���I�={C�O�s^?��}���?yKç'c�'sqH�`E�xp��������:!@I�>}@�n�@��@�: @l��?�٧]/ ���%�n�������=�=D���n/� ��@��oA�&{C/� @�U�/� �+J8���
H��>��=�3H��_�/ �F�6�G���E�A5F�ğ�E���/� ���fG��E���+E��E�X�?� >\�G��ZE�M�F?�lD�
`8? /�?n?�?�?�?�?�? �?O�?OIO4OmOXO �O|O�O�O�O�O�O_ �O3__W_B_{_f_x_ �_�_�_�_�_�_oo -oSo>owobo�o�o�o �o�o�o�o=( aL�p���� ���'��K�6�H� ��l�����ɏ���؏ ��#��G�2�k�V���@z�������韤"(�!�4�ퟦ���<�֕3�ϩ� ��!4 �{:�L��!��0+#f�x�Z��jb����1E����|�������쯠"��F�4���P޲Px�����������׿¿��湿����A� ,�Q�w�bϞ"$zό� �ϰ�����ߴ���@�.�d�R�ej�tߪߘ�0��������)�����.��R�@�v��  �2 H�6�&HY�����\��&B#L#B�  A� @'�����"�4�F�W���߁�������������$�� �� q�� ��%
 ��3EWi{ ���������* ��b�����4�$PAR�AM_MENU �?����  DE�FPULSE�+�	WAITTMO{UT�RCV�� SHELL�_WRK.$CU�R_STYL��OPT���P�TB��C�R_DECSN�i�<, 6/H/Z/�/~/�/�/�/ �/�/�/?? ?2?[?�VSSREL_IOD  �����j5�USE_PROG %e%W?�?k3CCR�|2��m�7�_HOST !Fe!�4O�:T���?-C�?A/CiO�;_TIME�|6�5�VGDEBUG�z0ek3GINP_�FLMSK�O�IT�R�O�GPGA�@ 2�Lp� [CH�O�H�TYPEbn� V?P?�_�_�_�_�_�_ �_oo?o:oLo^o�o �o�o�o�o�o�o�o $6_Zl~� �������7���EWORD ?	�e
 	RS��@�PNS���s�JO!�TyEP@}�COL�h3���3WL�0 ��՜
���5d�ATR�ACECTL 1��o .v�s ������|&���DT Q����S��D � �h�t��h� `�r��� ��	 ��$P������ğ ֟�����0�B�T�����j��r��������������j��r��R�� ���ޯ ���&�8�J�\�n�*�������Ȱk�U�r�����������Ȱܴܴ	ܴ
ܴ��޿���&� 8�J�\�nπ�Z���� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�X�j�|���� ����������0�B� T�f�x���\������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_���_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����_� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��� ����&8 J\n����� ���/"/4/F/X)��$PGTRACELEN  W!�  ���V �l&_UP ������!̣ �!� l!_C�FG ��%T�#V!� ��${#��/�(�-  ���%�"DEFSPD� ��,U!~ ��l IN� TRL' ��-�!8�%C1�PE_CONFI�� ��%��!�$�)l LID�#��-	�9LLB� 1�~7 ���$B� � B4�3�& ��5JOE�/ <o< T!?�1K PO1OHOjO�O~O�O�O �O�O_�O�O_L_2_T_�_�ZB�_�_�_ �_3O�_"oo'oXo�9�GRP 1��<�W!@�  �[��V!A?x�D� P�DV�C�2�� o�V d`,D�i�i�1�0��00Wo)O�1�n´(s
�kB+pRq2.h�R�V!>'oY>�a����~� �=N�=R� �3��0�i�T���x�����Տ������ G Dz0�9�V 
 � a��q���������ߟ ʟ��'��$�]�H�Ё�l�����)W!
�V7.10bet�a1�$ܠB�(�A�\)A��G��aޡ>�������ޡA�����ffޢ���A�p�AaG��Q�Q@�(��` ��K�]�o����#Apأ�r�0����Ϳ߿ ڢU!��}���v�$���H�2ϝ:KNOW_M  �%�&�4�SV ��9��5N����� f�9�$�6�o��"�m�3�Mvc���} ��	��"V ����T���Pܽ����פ�@1ߠ�`��(�wP�1MRvcĥ�T~�D��u������OADBANF�WD�ϡ3STva1� 1ś)��4 �5�����&��� � Q�D�V�h��������� ������
O.@ �dv�������2�����V �<%�w`3!3E���4bt����5 ������6//,/>/��7[/m//�/���8�/�/�/�/��M�A���d3�'O�VLD  ;��ߊ���PARNUM  ��?�?��SCHS9 a5
��7�1�9��
EUPD�?�5uTO�%_CM�P_��V0����'���lDER_CHKzE����ҎFwOƉKRSg���pa_M�O���H_�O�%_R�ES_G���;
 8��oi_\_�_�_�_�_ �_�_�_o�_/o"oSo Fo9?+U6\F_xo +Ua�o�o�o-S��o �o�o-S 27-S Z Rqv-S� ����-S 0���-RV� 1������@�`z$�BTHR_�INRg�X1����d�c�MASSp� Z愇MNo���MON�_QUEUE �������@���$N�q@U�AN��ۈ�E�ND��_�EXE ��6@BE���OPTIO��[���PROGRAM %Պ%�.��?~�TASK_IU4�g�OCFG ��Տ�?ɟ��DATA:����@�@M� 2 �f� (���������@c��΢֯�����ɣ  @6�>�P�b�t������INFO���I�� 䄽�ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/ߊ�4�����I� di��~�@DIT ����߬���WERFL�A�V���RGADJ� Ή�A�  ��?�@�w����� ���W��?�r��z��@<@�9���%?h���dm�C��2�%糲	H�lR7�U�2�?G�A �w�t$��*��=/�� **:���@�������5,�'�����1��1W�9�Q� ���/�A�o�e�w��� ����������] G=O�s��� �5��'� K]���/�� ���y/#/5/c/Y/ k/�/�/�/�/�/�/Q? �/?;?1?C?�?g?y? �?�?�?)O�?�?O	O O�O?OQOOuO�O_ �O�O�O�O�Om__)_ W_M___�_�_�_�_�_ �_Eo�_o/o%o7o�o@[omo�o�o�oN�	� <��*cNt�����Q�M���PR�EF �%������
��IORIT�Y��܆���MPDCSP�����C�U��|����ODUCT�������OG��_TG��钍ڂ��HIBIT_DO�A���TOENT �1Ӊ� (!?AF_INEm� �~+�!tcp+�>S�!udB�{�?!icmj�q�ւ�XY�ԉ����)� ��ߟ����ٟ���	�F�-� j�Q�c�����į���@�����B�T�*����%���V����>VӰ�f��/�	��������~��A~G�,  ���o�D�V�h�z��պ��Z뿺������ϻ��i�ENHANCOE �u�s�A��Ad�P�7�~����������PORT_WNUMn�������_CARTR�EP�Ĝ�SKS�TAm��SLGS6��ě�G�T��Unothin�gX�5�G�Y��{��T?EMP ڑ�e���e�_a_seiban����� ����"��F�1�j�U� ��y����������� ��0@fQ�u �������, P;t_��� ����//:/%/�^/I/[/�//�/q�VOERSIL���� � disab�lej�m�SAVE� ۑ�	26�70H755�(�/E?!@�G?Y?|�}?C 	�8w��o�;�?��e�?O"O4OFOTJA�<|?�O��5_��W 1�ě20�@�r�e�O�O�g�pUR�GE�B掘�WAFP�p����W��3T�ѯ�WRUP_�DELAY ����&UR_HOT �%!vz�?߳_DUR_NORMAL�X𙂢_�_�WSEMI��_�_;o�qQSKI%P�C�|��Cx�/�o �/�o�o�o�m}�o's �o!3EiW� ��w����� /��S�A�c������� s�я������ߏ� O�=�s�����]������˟���SRBT�IF4T��RCVT�MOU������/�DCR�C�^i� ЗaB.&��B���B'��w@�qy@��)ݹ4�m�,����e�p]2�?)���9��o�ݯ�o<2�!<"�7�<L��<`�N<D��<�A�ɫ0�ׯ@�Q�@� u���������Ͽ�����)�;�o�RDI�O_TYPE  ��M1�G�ED�T_CFG ��6KbBHSE��Xa�2�� �� ������.� �үD�/� h�S��ϙ�(o���o�� ӟ�����;�)�_�M� ��m�ߴ�9�{����� ���%��5�7�I�� �������a������� !E3i����� a�]��� A/e���mG ���/�+//O/ qv/�/G/�/C/�/�/ �/�/�/'??K?m/r? �/S?�?�?�?�?�?�? O�?!OW?}?nO;���?INT 2�Y��=�_�G;� �O�K��+��OX�f�0  _[3O6_'OF_H_Z_ �_~_�_�_�_�_�_o �_2oo*ohoVo�ozo �o�o�o�o�o
�o. @&dR�v�� ������<�"��`�N���!�EFPO�S1 1�d�  x\O҉���O ����+�ŏ׏�r� ]���1���U�ޟy�۟ ���8�ӟ\������� -�?�y�گů����"� ��F��C�|����;� Ŀ_���������B� -�f�ϊ�%Ϯ�Iϫ� ���ߣ�,���P�b� ���Iߪߕ���i��� �����L���p�� ��/����e�w��� ��6���Z���~��{� ��O���s����� 2 ����ze�9� ]����@� d���5G�� �/�*/�N/�K/ �//�/C/�/g/�/? �/�/�/J?5?n?	?�? -?�?Q?�?�?�?O�? 4O�?XOjOOOQO�O �O�OqO�O�O_�O_ T_�Ox__�_7_�_�_ m__�_oo>o�_bo��_�o!o�o�oUc��2 1崏^opo�o( LRop�/� �e����6�� ��/���{���O�؏ s�������2�͏V�� z����9�K�]����� ����@�۟d���a� ��5���Y��}���� ��ů��`�K������ C�̿g�ɿϝ�&��� J��n�	��-�g��� ���χ�߫�4���1� j�ߎ�)߲�M���q� �ߕ���0��T���x� ��7����m���� ���>�������7��� ����W���{��� :��^����A Se� �$�H �li�=�a ��/���/h/ S/�/'/�/K/�/o/�/ 
?�/.?�/R?�/v?? #?5?o?�?�?�?�?O �?<O�?9OrOO�O1O�OUO�O�o�d3 1��o�O�O�OU_@_y_ O�_8_�_\_�_�_�_ o�_?o�_co�_o"o \o�o�o�o|o�o) �o&_�o��B �fx��%��I� �m����,���Ǐb� 돆����3�Ώ��� ,���x���L�՟p��� ����/�ʟS��w�� ��6�H�Z������� ��=�دa���^���2� ��V�߿z�Ϟ���¿ ��]�Hρ�ϥ�@��� d����Ϛ�#߾�G��� k���*�d��߰��� ����1���.�g�� ��&��J���n��� ��-��Q���u���� 4�����j������� ;������4��� T�x��7� [��>Pb ���!/�E/�i/ /f/�/:/�/^/�/�/x?�OT4 1�_ �/�/?�?m?�?�/�? e?�?�?�?$O�?HO�? lOO�O+O=OOO�O�O �O_�O2_�OV_�OS_ �_'_�_K_�_o_�_�_ �_�_�_Ro=ovoo�o 5o�oYo�o�o�o�o <�o`�oY� ��y��&��#� \�������?�ȏc� u�����"��F��j� ���)���ğ_�蟃� ���0�˟ݟ�)��� u���I�үm������ ,�ǯP��t����3� E�W����ݿϱ�:� տ^���[ϔ�/ϸ�S� ��w� ߛϭϿ���Z� E�~�ߢ�=���a��� �ߗ� ��D���h�� �'�a�������
� ��.���+�d����#� ��G���k�}�����* N��r�1� �g���8?045 1�;?�� 1������/ �/Q/�u//�/4/ �/X/j/|/�/??;? �/_?�/�??�?�?T? �?x?O�?%O�?�?�? OOjO�O>O�ObO�O �O�O!_�OE_�Oi__ �_(_:_L_�_�_�_o �_/o�_So�_Po�o$o �oHo�olo�o�o�o�o �oO:s�2� V�����9�� ]��
��V�����ۏ v�����#��� �Y�� }����<�ş`�r��� ���
�C�ޟg���� &�����\�寀�	��� -�ȯگ�&���r��� F�Ͽj�󿎿�)�Ŀ M��q�ϕ�0�B�T� ������߮�7���[� ��Xߑ�,ߵ�P���t� �ߘߪ߼���W�B�{� ��:���^���������A���e�K]6 1�h�$�^��� �� �$��H��E ~�=�a�� ���D/h� '�K���
/� ./�R/��/K/�/ �/�/k/�/�/?�/? N?�/r??�?1?�?U? g?y?�?O�?8O�?\O �?�OO}O�OQO�OuO �O�O"_�O�O�O_|_ g_�_;_�___�_�_�_ o�_Bo�_foo�o%o 7oIo�o�o�o�o, �oP�oM�!�E �i�����L� 7�p����/���S��� ����6�яZ��� ��S�����؟s��� �� ����V��z�� ��9�¯]�o������ �@�ۯd�����#��� ��Y��}�ϡ�*�ſ ׿�#τ�oϨ�C��� g��ϋ���&���J����n�	ߒ�x���7 1��?�Qߋ�	���-� 3�Q���u��r��F� ��j����������� �q�\���0���T��� x�����7��[�� ,>x��� �!�E�B{ �:�^���� �A/,/e/ /�/$/�/ H/�/�/~/?�/+?�/ O?�/�/?H?�?�?�? h?�?�?O�?OKO�? oO
O�O.O�OROdOvO �O_�O5_�OY_�O}_ _z_�_N_�_r_�_�_ o�_�_�_oyodo�o 8o�o\o�o�o�o�o ?�oc�o�"4F �����)��M� �J������B�ˏf� ������I�4�m� ���,���P���럆� ���3�ΟW���� P�����կp������ ���S��w����6�x���߷�8 1��� l�~���6�!�Z�`�~� Ϣ�=ϟ���s��ϗ�  ߻�D������=ߞ� ����]��߁�
��� @���d��߈�#��G� Y�k�����*���N� ��r��o���C���g� ����������n Y�-�Q�u� �4�X�| );u����/ �B/�?/x//�/7/ �/[/�//�/�/�/>? )?b?�/�?!?�?E?�? �?{?O�?(O�?LO�? �?OEO�O�O�OeO�O �O_�O_H_�Ol__ �_+_�_O_a_s_�_o �_2o�_Vo�_zoowo �oKo�ooo�o�o�o �o�ova�5� Y�}���<�� `�����1�C�}�ޏ ɏ���&���J��G� �����?�ȟc��ҿ��MASK 1���0�>��XNO  �=�C��MOTE  _� � ��_CFG �휭��PL_RANG�������٦OWER ������SM_�DRYPRG �%��%��I��T?ART �	�W�UME_PRO&��8����_EXEC_ENB  ��=��GSPD��ΰvָ�TDB���RM��I_A�IRPUR� p��m�p��MT_��T�����OBOT�_ISOLC]���l�̥ȥ��NAM/E ������OB_ORD_N_UM ?	�i��H755 � ��@�R�d��P�C_TIMEOU�T� x�S23�2��1�`�� �LTEACH PENDAN��X��С��������Mainte�nance CoKns������"�����No Use �����@�R�d�v�����NPOf���С�����CH�_L�����	����!UD1�:1���R�VAI�L!ц�������S�PACE1 2�`�
��ХЩ�巓ΦТ�m����< ���?� Y�Y���KlC� |���������% <�QrY`�d� �����Y) /@/�U/v/]/�/� �����//7/-? �/Q?r?�?k?�/�/�/ �/�/�??3?)OJO	O _O�OgO�O�?�?�?�? �?OOAO7__[_|_ �_e_�O�O�O�O�O�_ _=_3oToou_�oqo �o�_�_�_�_�oo)o /Moe�]o�o �o�o�o�%G=� ^����{����� ����!�S�9����@o���g������2��� ��ݏ���� %�W�Z���:�������Ưǟ3ڟ����"� ԯF�x�{���[���ҿ����4����1� C���g������|��������	�5�.�@� R�d�߈ϺϽ�ߝ� �����)�*�6=�O� a�s߅�7������$�@���5��J�K�7^� p����X��������E���5V-kl�8 ���������y��  f VwN���G �� t�ń
� �  �//1/C/U/ g/y/���-���/m�/ȁd0�/2? D?V?h?z?�?�?�/�/ �.�:�?�;O??�? ZOlO~O�O�O�O�?�? �?�?O_5_(O:O�O z_�_�_�_�_�_�O�Op�O _"_4o `� @Ȁme�/{oW__Y�a�UDo�o�o�_ �j�o�o1CaI ��gq���� ���Q�c���7�i� ����������Տ�ُ��\
�ol��A���*SYSTEM*��V9.1018�5 ��12/11�/2019 A� �� ��r�ӓS�R_T   �� $ĐENB_�TYP   �$RUNNER�_AXS� $H�AND_LNGT�H�`�THIC=K��FLIPґ�`�$INTFER�ENCE��IF'_CH��I֑$�=9�INDXD�Đ�G1POS  � W�N�`�ANuG`�x�_JF���PRM`� 	�RV_DATAƑ�  $��E�TIME  ��$�VALU����G�RP_  � ��A  2� �SCő�	� �$ITP�_�� $NU�MڠOUِ	�TO�T�
�DSP!�J�OGLIM� $�FINE_PCN�T@�CO��$�MAX�TASK�@�KEPT_MI�R=�]�PREMT�q�}�APLD���_EX������t�@���PG��BRKHGOLD�!��I_��  ڲ@���P�_MADE�w�B�SOC�MOTN��DUMMY16�3�SV_COD�E_OPM�SFSPD_OVRD���R�LDL�O�OR�Z�TPӐLE[�F�!�[�:�OV=�SF��ᐓ�T�F��A�a��UFRA��TOO�L@�LCHDLY>W�RECOVK�퐆:�WSs�:��=�R�OM��I�_�ڐ� @��S��NVE�RT�OFS;�CǠD�FWDt���p���ENAB��7�T�R��`���E_F�DO��MB_CM����B-�BL_M�i�]��Ҫ�2S�VS{TAA�$UP��d���G�׸�AM��`��а��%� �_M���A�AM�A�1�T$SCA0�,�D�7��HBK���L�IO�?�[�IQ�$PPAO�{�`��s���s�1�DVC_DB ��F����쑼��A�"��1��%���3��+�/ATIO� �h��K�U��/�/�P�ABF�T֒E�G�Ԛ��ؼE�:�_AUX�S�UBCPU�G�S�IN_7Ў���P�18������FLA��ݑHW_C1���j�|����$ATR����$UNIT�|����ATTRI����G�CYCLC�N�ECA!�FLT�R_2_FIR�T�ARTUP_CN�`Ӷ�SIGNO�L�PS�2�1�_SCT6z�F_��F_��t���FSF����CH�A��[���O��RSD/���/�P��s�;_T��PRO�|ӎp�EMP�=��T����ܐ���'D�IAG�RAIL�AC��p�M�LOh��'�4�PS-�b@� i�+�%�PR��SB�  �Cް� 	$�FU�NC���RINS_TB���=�o�#RA��`�7��8a�E��WARq�8��BLCUR�$A0+	((DA��G(#%LD=�?�h��o#��to#TI���%�ܐ$CE_RIA_SWA�+AF��P^��#�6�%T2\CK��C�MOI���DF_�LE�_�PD�"L�M��FA�HRD�YO��E�RGt H�� z���O 5MUL�SE� ���0���$JW�Jrǂ�F�AN_ALMLV��Î1WRN�5HA#RDאO�_O,� :�2�1STO�ƵY_���AU��R�<(���_SBR���5�.�J���CMPINFڐ��-De!n8CREG@�NV0�l�$�۱DAL_N��FL����$M  2��7%�ܐ�8�E�CM-�N0�Y������G���SP$�R�$Y��Z�����ۡ��� ����EG!`
�?�
QAR�0�'�20�U3 AXE$�ROBn!�RED!�WR�2߱_i]�SYܰDQtᰋVS�WWRI�V��STR �)��
f�E��Ġ&To�1"�B�P1��V5c��OTOHAĠ�ARY�b]�ΡR��FI��h�$LI�NK�!��3a$E�XT_�S1�%U6��[aXYZ�2ej7NsfOFF9�2bZbJNh`B���d0�����cFI �g��A�7Ĩ9�_J L�¢d�?ch��0�T�[-8�US��B	qL22ArC7 ��DUO�$V]9pTUR�0X�#�zu!a(BX�P,�)wFL[`��@�P�p|e�Y�30�G� 1JĠKF�M�'�3���s�����a�ORQ .���x��s��m��� �H��,�_A]�OVEd���Mh l��C ~��C~��B}��0{�B� |���{�~��h� �� e�u�����l�v�e���`��C���.�ERK�
�	tEЪ��E�	A�ܐ�e� gN!K�N!AX�¢N! ���4b��0��Z1�� o��`��r`���`��:p��qp��1�p��:0 ��:0��:0Ǚ:0י:0 �:0��:0�:0�:0x'�D�8�DEBU��$��3(�N�VbCABNL�t�^�VA��� 
����+� ��7�0�7�o7�a7� ra7��a7�:q7�qq�$pFp�"ۂ�cLAB�bq)�����GRO: 4)r�<*�B_,� �Tm��`�0��*���1�AND�pt�:� +�_e=��1Y� *��A��Pm�!|�- ^`NT8�0ӟ�VELل���L���SERV9E���@ $�`�mA]!��PO@� � ��`���@���!�@  $�TRQ�r
 �tR
���"2�q I?_ 	 l���N[ERR�boI,�8��لr�TOQلրALHP���R�� G��i%Ha�����REP  
 ,��#�=��݁RA�� 2	 d��s��@���7 �@$r�l� ��z$ �OC?!��  d�C�OUNT�Q� ��SFZN_CFG�	� 4��aF3T ������ܣq ��L�Q�^�C �(�M���g2��Ճ{����F!A� 䅻&��XdP�� ����SQ��G�dQ9PB��@HEL}@Y� 5pB�_BAS��RSR`F�^SS��!M�1��M�2p�3p�4�p�5p�6p�7p�8��@�ROO�p��V f]`NL�ALsAB���FN�ACK�IN�Tg �CU�0E0�� 	_PUdq�2ZOU��P�aH-�֨ ��P��TPFWD_�KARw�iAf�RE���$0P/`U!w�QUE`I e�Up�r�0�1I�0�-�[`S��SF[aSEM3��A�0�A��STYSO� 	�DI�}�܄��!_TMuCMA�NRQL[`END��t$KEYSWITCH^s.��HEUpBEATM6�PEPLEv������UrF�sS~3DO_HOM� �O�1 EFA�PR��a�vQ�P�EC�Ox01c���OV_Mr<� � IOCMGt��A��B.�HK�A# DXabG��U^ҹ�MP�W�WsFORCfCWAR 2��.��OMP  @���c�0U�SP3P1(�&�@�$3�&4���*�O� L�"��aHOUNLO9 \�4�ED�1  �S�NPX_ASZ�; 0�@ADD���$SIZfA$�VA���MULTKIP��.3� A�! � $H	�/0��`BRS}�ϱC<rТ6FRIFu��aS� �)��0NFOODBU�P~��5�30�9�ƽAfIA�!$V��y�x�R�SN��@� � L0��TE��s8�:sSGLZATAb�p&o�sC᳍P[@OSTMT�q�CPP�VBWe�\DSHO�W�Ev�BAN�@TP�`�wqs8��s8��r���V7�_G�� :p$PCD �7���kFB�!PXSP� �A U�ADP���� �W�A00^�ZR� bW� bW� �bW� bW5`Y6`Y7�`Y8`Y9`YA`YB�`Y� bW��cV�@bWF `X7�$hlY(@$h�Y@@T$h�Y1�Y1�Y1�YU1�Y1�Y1�Y1�YU1i1i1"i2_YU2lY2yY2�Y2�YU2�Y2�Y2�Y2�YU2�Y2�Y2�Y2�YU2i2i2"i3_Y��p�xyY3�Y3�Y3��Y3�Y3�Y3�Y3��Y3�Y3�Y3�Y3�i3i3"i4_Y4�lY4yY4�Y4�Y4��Y4�Y4�Y4�Y4��Y4�Y4�Y4�Y4�i4i4"i5_Y5�lY5yY5�Y5�Y5��Y5�Y5�Y5�Y5��Y5�Y5�Y5�Y5�i5i5"i6_Y6�lY6yY6�Y6�Y6��Y6�Y6�Y6�Y6��Y6�Y6�Y6�Y6�i6i6"i7_Y7�lY7yY7�Y7�Y7��Y7�Y7�Y7�Y7��Y7�Y7�Y7�Y7�i7i7"d�VPz�U� ��߰e�
�A�2�� �x #�R�@  ��M��R9� ��Q_+�R����(�~ J��S/�C�D�^��_U�0i�C"YSL|���� � L5 Bj��4A7�D����&RVALUj�% x�1���F��ID_L��3��HI��I�"$FILE_L!�ic$�� ��SA�� h	�M�E_BLCK�Z�uAc�D_CPUs�M0sـA0u�$�6ԁ¯GR�  � PaW-����0��LA�A�S�������RUN_FLG���� ���v�!���!���H�F ��C�������T2x_LI�"�  ��G_O��� P_EDI0�"Y���c�k�9���nє0�!�TBC=2LT �Q@ 0�(0�!c�FT���.	TDC�A4z����M�������THD�0�!�#�$�R��<0e ERVE�F�	F�5A�� �  X -$q�LEN�~�	q�) cRA� 2��W_?�Ҡ�1q��2��MO$k�5S�0 I. Z�`����q���DE��1LACE,":�CqC3Z¶_MA20p>>TCVEfTXg
�|
8R�Q�QJAUM���J>JP)�}�2��@�BP	0JKV�K�A.)A.5A#J��AF2JJ:JJBAAL2h:h�bAAf5#� N1���XB G�L��_l�A�0IB��CF62�! `	�GROUP��vA�2$QN��C�3~�REQUIR1��0EBU�3m��$T 2 *!n�&8��50��" \� ��oAPPR  CLG��
$t�Ng(CLOD��w)S��)
��.u6# ���M �C 8� 2�$_MGA� �CLPN��(� R �'B{RK�)NOLD�&�@RTMOb�:
=�%Jb�4Pj  :�  B  �  �  6rW57W5hA  ��>��$� "����A�7)A�3PATH�7�1�3�1���3� r/ #\�PSCA��� 7h"�!INp�UCh����0@C:PUM9H	Y���� @A��L��[J�0[Jq0[@PAYwLOA7J2L�OR_AN��CL���I�A�I�A�%R_F�2LSHR@��AL�O�D~A�G=C�G=CACRL_��-E P)G�D;H��G�$H��"NRFLEXj#:��J��% PT"��`��E�W��Z�BJp�& :}���  �W�T��< ������F1�QEeYg������(�bE2DV hz����`x}t ��m`�x��$�QT�w^qXF�� �d�h%.�x1C Ugktb�����C�kP�' ������	/���ATrf!� EL�`(�D�j#(J/ &* JE0gCTR)AmaTN���@�'HAND_V�BG�jQ���4( M$�pF2�&����SW�Y���&)� $$M�@�)!� �!�1�#p��E2��A���@�&��<��-A(�,���*A;A;G���+���*D;D;P2�0G��ݩST�'�49�N8DY�e  �&(�O��@r��G�Q�G��A�G�t`�5P _5h5q5z5�5�5�5�2:�J��* ��T��2 �a㵙!�A'SYMEZ� F!)K� L�A$O_B�X 5@HD2=4ĸ�ROdOvO�O�CJ�LR0�J����L�Id_V�ׁ�<�#!�V_UN���6�W��AJN�|�N� �LR�U_ԃ�]� $Y R03_E_���[TcS�   �T��HR���+���}P]"DI0#O#�gR�N�, g�V�I9�AV1SP�s`^�^�v`�P����`� - �� ɑME�aЫ�y���`�T�PT@��Հ�0����V ��������T���� $DUMMY}1q1$PS_p`�RF2`�0$��n�PFLA�YP����$GLB_T��1���]!�P�`q�}�. XT '�1�ST�* SBR��0M21_V�T�$SV_ER�@O���w��CLK�w�A��`OS� �GL�E�W�/ 4���+$YX�ZX�W����AœAz�9B肼�U.��0 �pN����$GI��}$�� /�P������1 L���}�$F��ENEA�R�`NwcFd	�`T�ANCwb����JOG&`H0 2�2�$JOINT��"��1��MSET.�3  EJ�a��S���1��4�� n`U�a?��* LOCK_F�O�@Б�BGLV�t�GLTEST�_XMj �EMPĠ �r2I�� $1U�P��9`20* ��BX1#̐� X/y��CE�&y $K�AR$qM%�TPD�RA���VECX`�� IUX2]{HE TOOL9c��V8dRE�IS�3�U�6z1m`AC)H� / 3�O@��j��3g�% SIZ"�  @$RAI�L_BOXE�ޜ�ROBO)?�~��HOWWARVQxH!��!ROLM� n%ԁ$"�6 a`�0�O_F�!��HOTML5�)AͲ��!�15��R
�O�R6�"1`�� o 
��OU�'7 d��T/`�J�|$�� $PIP*N�p�6"!`X� ~�PCORDED� �
@� a XT*0)� � �O`� 8 7D 0�OB|�N� � �7v1��/�v2��P�wSYSv1ADRO�� ��TCH� 79 ,�pEN	�QA_�4݁@����VWVA|�:� � ����P�REV_RT���$EDIT(FVSHWR�c�G@�bJ���D��O�^D~W�$HEAD��h��x@��0CKE����CPSPD�FJKMP�0L�iPR�`F;�;~0{Q�6I35SO�C��NE�P����TICK9c��M��Qu�CHNY��< @�0�AᅗA_�GP&V-&�PSTY��2!LOK� ��D"R�P= t 5
#@G�5%$Au=c�SE�!$D� 9`���M��P&�&V�SQU�,e��TGERC��ʱv�S�>  o���p��q�``O����{`�IZ����P�R\0�Db�A0PU�;�Te_DOi�0XuS� K�AXIs`�#]UR��cP� O P�6���_��2�ET�bP�0	��rPF	�sPA�����9'[) ��S=R��?l�P� !���/u�Ay�/u*� /s8�/sH�uuj�uuz� uu���u�}���u�|���yC
��}C�}�ϕϸ�Ϲ�-SSC3� o@ h��DS4P̗��SPJࡅAT�x� �UaP�B��A_DDRES�B3@�SHIF�O_2+CHO��1IR����TUR�I�� }A�"CUSTO�d*�V�I>�B�2���8c�
2
ՒV81da~�C \a�8A�rPC�a�P��C���b�bR�6���T�XSCREEx2Dz��QTINA���# Ӕ) � Q_��ٰE T�A��8b �1��n� ��a�2�b�/@RROS�~ �0�@��o� ��UE��DF ���1
�S���1RSMPwgU`e0�P抡�S_�󀪦=Ú���ȧ=õaCx���� 2E� UEմGD���D`WGMT��Lp��a�~�O�04�BB�L_ W��~�H ��rPJ�O��V�L�E�a�N �`�RI;GHj�BRD��ہOCKGR����Tf0|����WIDTH#�T@n�)!����UI� EY��}�I�
2� m VR6 @aB�ACKTQ�Ũ���FOS1�LAB�_q?(��I ��$URT!E��I_���H@� J 8���~ _wA�h�R����s(��o0U�O��~�KP����U�v���Ry!LUM8�ØfՀERV!1��RްPh �L���`�GEI�O�`l2�@LIP��bE�Pf�)%�@v�3؆�3�  2�50�60�70�8��R��?`h ���� !�Sv�PKݱUSR��OM <a���U�(�FO�PR�I�am  ���TR�IP2!m�UN+DO;�N �P �ye`!xe@�O�`�P� Oc���CaG �PT� T��^�O	S��s�R�`F�J���Z�P��������6TA%CJ�U�Z�Q���pã�5UJ�OFF(�[�R_���O)� G1P���;�Q��GU�1P:��"V�Q�`��SUB6R���'SRT��tSR}̞ #cOR ��RA�U(p��T���7��_�&@�DT |1p�8O�WNM��4$SRCQ�Ҡ�PD(&r�MPFIMTl��`ESPPab����eA����i���A@
�U M`��WO[p�4an�PCOP��$�`�O�_- b�1�WA3@CF�� Z����@l"+� V~�SHADOW�`���_UNSCAp��ʴDGD!��1EGAC�8���VCWp`
�Wǔ ,"w1�S$NER�c�Q#+�yC0cDRIV6f�a_V/P��@m �D��MY_UBY ��kyV��UR��P�beA�� "P_�MT"LZkBM]��$�@DEY�3EXX7�^��MU�@X]��V$��US���`�_�R�����
�R��QG>�pPACIN�A�PRG�$�"�"���"ң�RE}�遚��c�H�"@X �� G�P��� R�IR��@Y��?�dӱ��	�qaREb#�SW� _A�!e�$W#B`O��ہA�^3�/rE��UeP�d��@�IHKjRZ���v:�P&q[0%��3EA�P�7� j�^5۰IMwRCV
�[ ��UOvPMj�C��	�28��#�2REF6�F �6�1M0���c50���:�FAJFAKhE�6�?_  �:�H�;�pS��N'��aaQ�I�\ ��GR�ӵ`�м��POU4W�"Vk �W 5U�2��$0Ԑ��C`,�Y��U��2Q{�ՀULj�Zf_ CO~��[H EPNTZ�T��U���V�ђSQPL��U#�U���W���VIsA_���] �T��HD����$JO���6��$Z_�UPL�W�Z|pW�!e�QPSp�0�_LI��$EPEQ��k�@a�QǑ΁��΀K�P|]m�^� 0����a� ��CACHLO:A�d�aI �ih��� 1CI`MI惉FHa�eT�p�f�K$�HOj��`COMM���Ot�wW�Ӳ�S&�T7 VPx�"@�mr_SIZwtZ� rx!asw����MP�zFAI!`G��4�`AD�y�McRET�r|wGP���> & �ASYNB{UF�VRTD��%�|q��OL�D_���A�W��PC��T�U7#�`Q{0	�EC;CU�(VEM� �e<���gVIRC�q9��!���%�_DELA`�#&Q���AG5�RK!XYZ̠��K!�W1��8A��򱦀TN8"IM߁8�������eGRABB��YRb"C�e�_e���LAS��r1�a_GE�e`u�&��;����T/S&N` ���%I����"ņ�BGf�V5��PK� ǆ�aWKGI��N#�`2F�@��`�qq�a+�aS��p�fN:��PLEX��b�����;��Nq��I? �-|�� |�.$�3����- �"c��b�t�Ŀ��.}�ORD���1�иw�RN�d $MPTIT� �C��F��VSF����e a -�[�QK UR�6�SM!�f+���AcDJ�N%�PZD>�gg DƨBaAL+`x�p�AbPERIs`���MSG_Q9��$}q�u����b��h�+�"�g�J`�3p�X�VR#�in�b�T_�OVRi��ZABC��j�";�s/@?
nda�Z]�#�k+�=$L�-B��aZMPCF��l�H���A����LN�Kc�
m����m $,q�0�įCMCM� C�C����p4P_A+A'$J����Dbq� ��� �� ����
D��F�UX���UXE]!f��	�]��]��oс�oё���FTFpsQӾ�r1��Zbŏn {�}�L�����YJ`D�� o�Y�R�pU�$H�EIGH�#"�?(�MP�.A\����Dp� � EX�$B�QPx �SHIF,�s��RVI`F��/B|�0�C`�dTF @{"�������WuD��_TRACE��V�A�9� PHER� q ,MP�)�;�	�$R�!p�� ����F�� S�6�S � F��  �S�x�2p������ s���r�����	���U�C�ADC����l6�R   d�� ZD �Qx0C���l�l0�| ʆ6�V��@ 2�F���� D��P�����	�	F� ,:$ZH~l� ������ // D/2/h/V/x/�/�/�/ �/�/�/
?�/??.? d?R?�?v?�?�?�?�? �?O�?*OONO<OrO `O�O�O�O�O�O�O�O __8_&_H_n_\_�_ �_�_�_�_�_�_�_�_ 4o"oXoFo|ojo�o�o�o�o�o�oF��$S�AF_DO_PULSC�G��k�$qp����|k���5qR� ��`��XP�+S�S�
������s��tq  ���������*�<�N�`�r�����]�  ��2��Dtqtqd�������rs�� @�������*�܉�� � 6���_ @J�T�Y J���������T D������� �)�;�M�_�q����� ����˯ݯ��~�����M�_�8$��sR�;��f����p���
�?t��Di��q>��  � ���� R�q|ulq���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e�@w�����S��G� ������0�B�T�f� x������������ ��"4FK��b0E�ҳD�ܽ��� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?��? �?�?�?�?�?�?	OO -O��QOcOuO�O�O�O �O�O�OLz��!_ 3_E_W_i_{_�_�_�_ �_�_�_�Yoo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������ø��Ǔ�6�H�Z� l�~�������Ə؏ꏀ��� �2�D�V�d�p#�m�����������i�	123�45678ݲh!B!ܺT
z1!���
��.� @�R�d�v�������"� ïկ�����/�A� S�e�w���������ѿ ������)�;�M�_� qσϕϧϹ������� ��%�7����m�� �ߣߵ���������� !�3�E�W�i�{��L� ������������/� A�S�e�w��������� ������+=O as������ �'9��]o �������� /#/5/G/Y/k/}/�/ N�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�/	OO-O?O QOcOuO�O�O�O�O�O��O�O__)_;_BS��]_o_�?�_�_�_�ԚCz  Bp��z   ��2��� } �X
~g�  	��R�2U_<oNo`oro�l��\�+o�o�o�o�o "4FXj|� �������� �oB�T�f�x������� ��ҏ�����,�>��P�b�t����������Qa�R<Ք �˕a  ��������#a#at�  �P#�;���`��$SCR_GR�P 1�*P��3� � ���R �U	 ����������Qԑ�U�������ٯǯ ��]ٰ`��C�,�����m��C����lL�R Mate 2�00iD 567�890!`LRM�|� 	LR2D� ���
123	4��Ц�d��hbճ���}�ݣ}��cDԑ����ѡ�	j�4�F�X�j�|τ����H���Ē� }���į������̦<��1��A���e��WV���Vh`,R��o  ���B��P!ư߮��Ԫ�A�P���  @�0�ժ�@������ ?4���H��P'��ڪ�F@ F�`Q�Y�P�}�h� ������������� ʩ�����J�5�G�Y�k�B�y�������� ����=(aL �p��o�
'�����W`�.4�=@4�>�1U4̧�@��n�PȄ@����ݣT_��A��������aĲ�1 
/1/C/Q*!!f(r/�/S/�P�#
b�/�/�/� ?�/�$?,4]�ECLVLw  �1�����>1L_DEFA�ULTF4������0Z3HO�TSTRf=�z2MIPOWERFE0��Ur5�4WFD�Og6 r5=2RV?ENT 1M1M1��3 L!DU�M_EIP,?H��j!AF_IN�Ef0+O3D!FT$OZN!O~O!�ϣO� �mO�O!RPC_MAIN�O�H��O_�CVIS��O�I�_b_!TMPUPPUY_IdQ_��_!
PMON_�PROXY�_Fe �_�_uR�_Mf�_Fo�!RDM_SR�VGoIg5o�o!�R���oHh�o�o!%
�@MoLi�o*�!RLSYNC�+Qy8v!gROS O�|�4e��!
CEwPMT'COM�Fk��{!	�rCONS��Gl�Z�!�rWOASRCaoFmI�v��!�rUSB��Hn���O�Uc� ��?�d�+���O���s��П87RVICE_�KL ?%�; �(%SVCPR#G1ן�	�2�$�"�3G�L��4o�t�"�5�����6��į�7�����/�*�	97�<���od�� ����9����a�ܿ �������,��ٯ T���|��)���� Q���6�z���6���� 6�ʿD�6��l�6�� ��6�Bϼ�6�j���6� ���6���4�6���\� ^�
�ܟ������� ��.������8�#�\� G���k����������� ����"F1X| g������ 	B-fQ�u �����/�,/ /P/;/t/�/q/�/�/ �/�/�/�/??(?L?�7?p?�_DEV ��9�UT�1:|?�0GRP �2
�5�0�bx� 	� 
 ,�0x?�?�2�?OO @O'O9OvO]O�O�O�O �O�O�O�O_*__N_ 5_r_�_�?�___�_�_ �_o�_&o8oo\oCo �ogoyo�o�o�o�o�o �o4�_)j!� u������� �B�)�f�x�_����� ��������M�,�� P�7�t�[�m�����Ο �����(��L�^� E���i������ܯ��  ����6��Z�l�S� ��w��������ѿ� ��2�D�+�hϿ�]Ϟ� U��ϩ��������� @�R�9�v�]ߚ߬ߓ� �߷�������*��N� `�G��k������ �����&�8��\�C� ����y���������C� ��4F-jQ� ������� B)fx_��� �����/,// P/7/t/�/m/�/�/�/ �/�/?�/(??!?^?.e3d �e6	L?�?��?�?�?�?�?OK%��O5O<C��� NA�1NE^OlGVO�OzO �O�O�O�I"O_JI�O 4_"_X_F_h_j_|_�_ �O�__�_o�_0oo ToBodo�_�_�o�_�o �o�o�o,P�o w�o@�<��� ��(�jO����� p�������܏ʏ �B� '�f���Z�H�~�l��� ����؟���>�ȟ2�  �V�D�z�h�����ů ׯ��������.��R� @�v�����ܯf�п�� ����*��Nϐ�u� ��>Ϩϖ��Ϻ����� ��&�h�Mߌ�߀�n� �ߒ��߶���.�T�%� d���X�F�|�j��� �����*�����.� T�B�x�f�������� ������*P> t�����d��� �&L�s� <������/ T9/K//$/�l/�/ �/�/�/�/,/?P/�/ D?2?T?V?h?�?�?�? ?�?(?�?O
O@O.O POROdO�O�?�O O�O �O�O__<_*_L_�O �O�_�Or_�_�_�_�_ oo8oz__o�_(o�o $o�o�o�o�o�oRo 7vo jX�|� ���*�N�B� 0�f�T���x������ �&�����>�,�b� P���ȏ����v���r� ����:�(�^����� ğN�����ȯʯܯ�  �6�x�]���&���~� ����Ŀƿؿ�P�5� t���h�Vό�zϰϞ� ���<��L���@�.� d�R߈�v߬������ �����<�*�`�N� ���߫���t������ ���8�&�\������ L������������� 4v�[��$�|� ����<!3� �T�x��� �8�,//</>/ P/�/t/�/��//�/ ?�/(??8?:?L?�? �/�?�/r?�?�? O�? $OO4O�?�?�O�?ZO �O�O�O�O�O�O _bO G_�O_z__�_�_�_ �_�_�_:_o^_�_Ro @ovodo�o�o�o�oo �o6o�o*N<r `���o��� �&��J�8�n���� ��^���Z�ȏ���"� �F���m���6����� ����ğ����`�E� ���x�f��������� ����8��\��P�>� t�b���������$��� 4�ο(��L�:�p�^� ��ֿ�������π��� $��H�6�l߮ϓ��� \��ߴ������� �� D��k��4����� ���������^�C��� �v�d����������� $�	������<r `������ � $&8n\� ������/�  /"/4/j/��/�Z/ �/�/�/�/?�/?r/ �/i?�/B?�?�?�?�? �?�?OJ?/On?�?bO �?rO�O�O�O�O�O"O _FO�O:_(_^_L_n_ �_�_�_�O�__�_o  o6o$oZoHojo�o�_ �o�_�o�o�o�o2  V�o}�FhB ���
��.�pU� ����v�������� Џ�H�-�l���`�N� ��r�������ޟ �� D�Ο8�&�\�J���n� ����ݯ������ 4�"�X�F�|������ l�ֿh�����0�� Tϖ�{Ϻ�DϮϜ��� �������,�n�Sߒ� ߆�tߪߘ��߼��� �F�+�j���^�L�� p����������� ���$�Z�H�~�l��� �����������  VDz�����j ����
R �y�B���� ��/Z�Q/�*/ �/r/�/�/�/�/�/2/ ?V/�/J?�/Z?�?n? �?�?�?
?�?.?�?"O OFO4OVO|OjO�O�? �OO�O�O�O__B_ 0_R_x_�O�_�Oh_�_ �_�_�_oo>o�_eo wo.oPo*o�o�o�o�o �oXo=|op^ ������0� T�H�6�l�Z�|�~� ��Ə��,��� �� D�2�h�V�x�Ώ�ş �������
�@�.� d�����ʟT���P�ί �����<�~�c��� ,���������ʿ�޿ �V�;�z��n�\ϒ� �϶Ϥ�����.��R� ��F�4�j�Xߎ�|߲� �����ߢ��ߞ��B� 0�f�T���߱���z� ���������>�,�b� �����R��������� ����:|�a��* �������B h9xlZ�~ ����>�2/ �B/h/V/�/z/�/� �//�/
?�/.??>? d?R?�?�/�?�/x?�? �?O�?*OO:O`O�? �O�?PO�O�O�O�O_ �O&_hOM____8__ �_�_�_�_�_�_@_%o�d_nQ�$SERV�_MAIL  �nUd`�JhOUT�PUTYh�oP@NdRV 2��V  g` (��Q4o�oNdSAVE�zlhiTOP10 �2�i d  j_ 2DVhz� ������
�� .�@�R�d�v������� ��Џ����*�<� N�`�r���������̟�ޟ����U�eYP��oKcFZN_CF�G �U�gc�d�a�eT�GRP� 2^��a ,�B   A��nQD�;� B��� � B4�cRB{21�fHELLW�C�U�f�`�ou�|��%RSR� �)�b�M���q����� ο��˿��(��L��7�pςϔ��  �a%�����Ϣ�����oP������S��Ǫ�2oPd��|��ɦHK 1׫ ߈߃ߕߧ� ����������%�7� `�[�m�������~ìOMM ׯ��ȢFTOV_E�NBYd�a�iHOW_REG_UI7��LbIMIOFWD�L����l�WAIT4���v���t`rX��d��TIMX�7����VAX`��>l�_UNIT3�v�iLCQ�TRYX���eN`MON_�ALIAS ?e��`heo�� ���
t��# �GYk}�:� �����/1/C/ U/g//�/�/�/�/l/ �/�/	??-?�/Q?c? u?�?�?D?�?�?�?�? O�?)O;OMO_OqOO �O�O�O�OvO�O__ %_7_�O[_m__�_�_ N_�_�_�_�_o�_3o EoWoioozo�o�o�o �o�o�o/A�o ew���X�� ����=�O�a�s� �������͏ߏ��� �'�9�K���o����� ����b�۟������ "�G�Y�k�}�(����� ůׯ鯔���1�C� U� �y���������l� ���	��ƿ?�Q�c� uχ�2ϫϽ������� ���)�;�M�_�
߃� �ߧ߹�d������� %���I�[�m���<� �����������!�3� E�W�i���������� n�����/��S�ew����$S�MON_DEFP�ROG &����� �&*SYSTEsM*�� 	��RECALL ?�}�	 ( �}�3xcopy f�r:\*.* v�irt:\tmp�back*=>1�92.168.1�.15:1666�8 PYk}�}4!a);MX����
xyzra?te 11 ����a/s/�/�!%61A/R@/R/�/�/? /�/�/�/a?s?�?�/ �/<?N?�?�?O?(? �?�?]OoO�O�?�?8O JO�O�O�OO$O�O�O Y_k_}_�O�O4_F_X_��_�_�_8"s:o�rderfil.dat/,�_�_hozo��o}/"mdb: ,/EoRQo�o�o�  3/�_�ogy�� /A�_��	�/� ��c�u����_B��_ P�����*_��Ώ _�q�������:�L�ݟ ���&���ʟ[�m� �����6�H�ٯ��� �"���Ưدi�{�� ��2���V������ ��,�Կe�wωϜ�D� @�R��������Ͼ� ��a�s߅ߘϪ�<�N� ������(ߺ���]� o��ߦ�8�J����� ���$����Y�k�}� ���4�F�X�������  o2o�o��gy��o 9�oT��	/� �Rcu��+= ����/*�N _/q/�/��C/��/ �/?&�J[?m? ?��5?��?�?�? /"/4/�?�?iO{OO��/;O�/VO�O�O_ ��$SNPX_A�SG 2����,Q� �P 0 '%?R[1]@J0_WY?�C%W_�_f_ �_�_�_�_�_�_o�_ 7oo,omoPowo�o�o �o�o�o�o�o3 W:L�p��� ���� �'�S�6� w�Z�l��������Ə ����=� �G�s�V� ��z���͟��ן�� '�
��]�@�g���v� �������Я��#�� G�*�<�}�`������� ׿��̿���C�&� g�J�\ϝπϧ��϶� ������-��7�c�F� ��j�|߽ߠ������� ����M�0�W��f� ������������� 7��,�m�P�w����� ����������3 W:L�p��� ��� 'S6 wZl����� /��=/ /G/s/V/ �/z/�/�/�/�/?�/ '?
??]?@?g?�?v? �?�?�?�?�?�?#OD�TPARAM �,U6Q ��	�'JP'D�@�'H~D�-PPO�FT_KB_CF�G  fC2USO�PIN_SIM  ,[sF�O�O�O�v@=@RVNORDY_DO  }E��ERQSTP_DSB�NsBU_aX�=@SR �I� � &�@TYL�E1a_�\�T�CT�OP_ON_ER�R_;B�QPTN ��E�P��C�RRING_P�RM�_0RVCNT?_GP 2�E�A�@x 	Q_Poh@`>owobo�olWVD%`�RP 1LI�@ �axI�g�o�o�o EBTfx��� ������,�>� P�b�t�������яΏ �����(�:�L�^� p���������ʟܟ�  ��$�6�]�Z�l�~� ������Ưد���#�  �2�D�V�h�z����� ��¿����
��.� @�R�d�vψϯϬϾ� ��������*�<�N� u�r߄ߖߨߺ����� ����;�8�J�\�n� ������������ �"�4�F�X�j�|��� ������������ 0BTf���� ����,S�Pbt����bP�RG_COUNT�F��R�ENB�o�M��D/_U�PD 1{[T  
�gBR/d/v/ �/�/�/�/�/�/�/? /?*?<?N?w?r?�?�? �?�?�?�?OOO&O OOJO\OnO�O�O�O�O �O�O�O�O'_"_4_F_ o_j_|_�_�_�_�_�_ �_�_ooGoBoTofo �o�o�o�o�o�o�o�o ,>gbt� �������� ?�:�L�^��������� Ϗʏ܏���$�6� _�Z�l�~�������Ɵ������_INF�O 1@%9& H�	 �c��N���r�?���@B�z=���t���	�@���>�!�vm��´�B������=�` @ߚ @���>��� >���� �C�/�CQ��Ch<C3����u��B������C�0B���Ã�G����9lw7�/���YSDEBUG��A ��d))Q�S�P_PASS��B?c�LOG u=�J!  �9���  �%!�UD1:\��<#���_MPC��@%H�#�@!̱A� @!~�SAV ��`�y���вC�׸�SV�TEM_T�IME 1���K  0  ���C������MEMBK  @%�%!����%�7�G�wX|& � @G���iߎߞ�b��߲����^� y�@ ����*�<�v�T�f�`x������ ��� ����
��.�@�R�d�v��e���������� ��(:L^p ������� ��SK�����@hRdX�� "�Q2sߣ�p�� �� �������%/7/I/[/O�u$� �u/�����/�/�/���/���?'?9?K?]?o?�$ s?�?���?�4^�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_�_)�T1SVGU�NSPDy� '�c��4P2MODE_LIM ��dg�0T2=P]Q���/UASK_OPTGIONX��g��Qw_DIr�ENB���5c��QBC2_GRP 2#c���_�"� C�c(\BCCFG !�[�~� o"Ekem`eo���o�o�o�o�o �o�o?*cN `������� ��;�&�_�J���n� ����ˏݏ�Ȍ�� ɏ*�<����r�]��� ����H�ڟԯ��� ��,��P�>�t�b��� ����ί������ :�(�J�p�^������� ��ܿʿ�� �6�� �J�\�zόϞ���� ���������.�@�� d�R߈�v߬ߚ߼߾� �����*��N�<�r� `����������� ��$�&�8�n�\��� HϪ���������|�" 2XF|��n ����� 0fT�x��� ��/�,//P/>/ t/b/�/�/�/�/�/�/ ��
??:?L?^?�/�? p?�?�?�?�?�? O�? $OOHO6OlOZO|O~O �O�O�O�O�O_�O2_  _B_h_V_�_z_�_�_ �_�_�_�_�_.ooRo ?jo|o�o�o�o<o�o �o�o<N`. �r������ �&��J�8�n�\��� ����ȏ���ڏ��� 4�"�D�F�X���|��� hoʟܟ������B� 0�R�x�f��������� �ү���,��<�>� P���t�����ο��� ��(��L�:�p�^� �ςϤϦϸ������ ȟ*�<�Z�l�~��Ϣ� �߲�������� ��� D�2�h�V��z��� ������
���.��R� @�b���v��������� ����N<r (ߊ����\��8&\Fz��$TBCSG_G�RP 2"F�  �z� 
 ?�   ��������@5//Y/k+~�$��d@ ��!?>z	 HBLk(z��&j$B$  C�`��/�(�/�/Cz�/�(=A�k(333?&ff?��i%�A��/m?80 k(c�͎6S5�0DHp?�=@�H0j%K1�5j$�1D"N!�?�?�?�? ;OJ�(I&�(nE�OLO ^O�O�O�O�O�O_ [��H:Q	V3.�00�	lr2d S	*\PTTy�k_*_ �Q�I 8�Pt]�_  �_�_,�[~J2�%�=Q�o�UCFG '�F� �"j��Lb�R"owh�wo�o�jO�o�o �o�o�o=(a L^������ ���9�$�]�H��� l�����ɏ��Ə��� #��G�Y��� d�v� ��2�����˟�ܟ�  �9�$�]�o�����N� ����ۯƯ��zf 6�BF�H�Z���~��� ��ؿƿ����2� � V�D�z�hϞόϮϰ� �������
�@�.�d� R�tߚ߈߾߬����� �����>�`�N�� r���������� &���6�8�J���n��� ������������" 24F|j��� ����B0 fT�x���� �/�,//P/>/`/ �/0�/�/�/l/�/�/ ???L?:?p?^?�? �?�?�?�?�?�?O O "OHOZOlO&O|O�O�O �O�O�O�O_�O_ _ 2_h_V_�_z_�_�_�_ �_�_
o�_.ooRo@o vodo�o�o�o�o�o�o �o*�/BT �������� �8�J�\��l����� ����ڏ����ʏ4� "�X�F�h���|����� ֟ğ���
���T� B�x�f���������Я �����>�,�b�P� r�t�����6Կ��� ��(��8�^�Lς�p� �ϔ������� ߾�$� �H�6�X�~ߐߢ�\� n��������� ��D� 2�T�z�h������ ��������
�@�.�d� R���v����������� ��*N`
�x ��F���� $J8n��P b����/"/4/ F/ /j/X/z/|/�/�/ �/�/�/?�/0??@? f?T?�?x?�?�?�?�? �?�?�?,OOPO>OtO bO�O�O�O�O�O�Ol �_._�O_L_^_�_ �_�_�_�_�_ oo$o 6o�_ZoHojolo~o�o �o�o�o�o�o2  VDfhz��� ����
�,�R�@� v�d���������ΏЏ ���<�*�`�N��� ��@_����ҟ|��� &��6�8�J���n��� ��ȯگ�����"���F�0�  l�p�� p���p��$T�BJOP_GRP� 2(8��  ?�p�i	����*���@���@�� 0�� � � � � �� �p� �@l���	 �BL�   �Cр D����<��E�A�Sʿ<�B$�����@��?�33C�*���8œ���� �2�T�����;��2�t��@/��?���zӌ��-�A�>�Ⱥ�� 0�����l�>�~�a߾s�;��pA�?��ff@&ff?G�ff�ϵ�8� ���L���}������:v,���?L~�}ѡ��DH��5�;�M�@�#33`�����>��|�<���8���`ự�	�D"���������`�r�|���"�9������g�v��x� �נ������������� 0(V�b������p�C�p�	���	V�3.0�	lr2d��*b��k��p{ E8�� EJ� E\�� En@ E��E��� E�� E��� E�� E��h E�H E��0 E� E}ϒ�� E��� E�x E��X F��D��  D�` E}�P E�U$�0�;�G�}R�^p Ek��u������(^�� E�����X 9�IR4! H%�
z�`/r"p�v#Ѭ߱/��ESTPARSI �d�����HR� AB_LE 1+��J %p��(�' �k)
�'�(�(o�w��'	�(
�(�(5p��(�(�(K!�#'RDI�/��?? (?:?L?^5�4O�?�;@�?�?O O2N�"S�?�� �:�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo�� �@�O��7�isO�O�O �OU?g?y?�?�?�8�"~pbNUM  8������x� �J K �"_CFG �,Y{s�@��IMEBF_TT�!pu��� �vVERI#��a�v�sR 1-��+ 8mp�dk�� ;��o  � ��,�>�P�b�t��� ������Ώ����� (�:���^�p������� ��ʟܟ� ��$�6� H�Z�l�~�������Ư د���� �2�{�V� h���������¿Կ濐��
��"�q_Sq�v@��u� MI_CH�AN�w �u u�DOBGLV���u�u��!x�ETHERA�D ?�%���v �������(x�oROUT�p!WJ�!*�H��SNM�ASK���s��255.��N�ߖߨ��N� OOLOFS�_DI� BŪ�O�RQCTRL !.�{>Cw/&�T�J� \�n��������� �����"�4�F�X�j��z��������#PE?_DETAI�����PGL_CONF�IG 4Yyiq���/cell/�$CID$/grp1��;M_q�9C�߮���� �,>Pbt� �����/� �:/L/^/p/�/�/#/ �/�/�/�/ ??�/6? H?Z?l?~?�??1?�?@�?�?�?O O�n}�? VOhOzO�O�O�Oq���O�M��?__1_C_ U_g_�?�_�_�_�_�_ �_t_	oo-o?oQoco uoo�o�o�o�o�o�o �o);M_q  �������� %�7�I�[�m����� ��Ǐُ�����!�3� E�W�i�{������ß ՟������/�A�S� e�w��������ѯ������ �U�ser View� )	}}1234?567890J�\� n���������5�	̿��0�2=���� π2�D�V�h�ǿٿ7�3 �����������o�1�߾4��j�|ߎߠ� ����#���߾5Y�� 0�B�T�f�x��ߙ�߾6���������,���M�߾7�������@������?�߾8u� :L^p������� lCamera;�1�@0BT2BE� ~��H�����//�  ��� f/x/�/�/�/�/g�/ �/?S/,?>?P?b?t?�?�����?�?�? �?OO,O�/PObOtO �?�O�O�O�O�O�O�? �7XىO>_P_b_t_�_ �_?O�_�_�_+_oo (o:oLo^o_�72+�_ �o�o�o�o�o�_* <N�or���� �so���a�(�:� L�^�p�������� ܏� ��$�6���7 t�͏��������ʟܟ �� ��$�o�H�Z�l� ~�����I��7(	9��  ��$�6�H��l�~� ��ۯ��ƿؿ������ǧ9��O�a�sυ� �ϩ�P������Ϙ�߀'�9�K�]�o߁�
	�0߼�������� ��:�L�^�߂�� �������ߕ�� � ��5�G�Y�k�}���6� ������"���1 CU���I+���� ������1C �gy����h �յ;X//1/C/U/ g/�/�/�/��/�/ �/	??-?��![�/ y?�?�?�?�?�?z/�? 	OOf??OQOcOuO�O �O@?��k0O�O�O	_ _-_?_�?c_u_�_�O �_�_�_�_�_o�O� �{�_Qocouo�o�o�o R_�o�o�o>o);�M_qm   i���������0�B�T�f�   v~������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~��������ƿؿj�  
`(�  �p( 	 ���B�0�f� Tϊ�xϚϜϮ���������,���� ��oq߃ߕ����� ������c`�=�O� a�߅�������� &���'�n�K�]�o� ��������������4� #5GYk���� ����� 1C�gy��� ����	/P-/?/ Q/�u/�/�/�/�/�/ /(/??)?p/M?_? q?�?�?�?�/�?�?�? 6?O%O7OIO[OmO�? �O�O�O�?�O�O�O_ !_3_zO�Oi_{_�_�O �_�_�_�_�_oR_/o AoSo�_wo�o�o�o�o �oo�o`o=O as���o�o�� �8�'�9�K�]�o� ��������ۏ��� �#�5�|�Y�k�}�ď ����şן���B�"�@ �*�<�N���$����+fr�h:\tpgl\�robots\lrm200id���_mate_��.xml
���Ưدꯀ��� �2�D�V�F���`���������Ϳ߿ ���'�9�K�b�\� �ϓϥϷ��������� �#�5�G�^�X�}ߏ� �߳����������� 1�C�Z�T�y���� ��������	��-�?� V�P�u����������� ����);R�L q������� %7NHm �������/�!/3/E.g��� �$�r�<< p� ?�E+�/E/�/ �/�/�/�/?�/?<? "?4?V?�?j?�?�?�?��?�?�?�?
O8OF���$TPGL_O�UTPUT 7|P�P� h tE�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o�o'otEh �=@23�45678901 Lo^opo�o�o�o�cF� Io�o�o�o/�o�3ew���Ez} �����'��� ]�o���������O�ŏ ����#�5�͏C�k� }�������K�]���� ��1�C�۟Q�y��� ������Y�ϯ��	�� -�?�ׯ�u������� ��Ͽg�ݿ��)�;� M��[σϕϧϹ��� c�u���%�7�I�[� ��iߑߣߵ�����q� ���!�3�E�W���HA}c!�������������@j/�.�p* ( 	 1oc�Q� ��u������������� ��)M;q_� ������ 7%GI[��?f�f &��-� #/5//Y/k/9j��/ �/H/�/�/�/�/?,? �/0?b?�/N?�?�?�? �?�?>?�?O�?OLO ^O8O�O�O�?|O�O�O vO __�O_H_�O�O ~_�_*_�_�_�_�_�_ ol_2oDo�_0ozoTo fo�o�o o�o�o�o�o .@dv�o^� �X����*�� �`�r���������� ޏ<�N��&���2�\� 6�H��������ڟt� Ɵ�"���F�X���@� ��(�z�į֯����� j���B�T��x���d� �����0���Ϣ�� >��*�tφ�俪ϼ� VϨ�������(�:���)WGL1.X�ML��o��$TP�OFF_LIM ������}�N_SV��  �����P_MOoN 8������2y�STRTCHK 9������VTCO�MPAT��6��VWVAR :�ݹY�� � �q������_D�EFPROG �%��%ZAD?15 ADR*����z�_DISPLA�Y���ޡ�INST�_MSK  ��� ��INUSE9R,���LCK5����QUICKMEN�Y���SCREx���7�tps�c��5����ҩ�_��ST*��RAC�E_CFG ;���Y���	z�
�?���HNL 2!<��`� ��L ^p������
���ITEM 2=�8 �%$12�34567890<1  =<)O<ai  !ow��3�z��A //w)/��v/� �/��/�/M/=/O/a/ {/�/�/�/U?{?�?�/ �??'?9?�?]?	O/O AO�?MO�?�?�?qO�O #O�O�OYO_}O�OX_ �Os_�O�_�__�_1_ �_og_'o�_7o]ooo �_{o�_	oo�o?o�o #�oG�o�o�oS k��;�_q :��U��y������ �%��I�	�m��?� ŏ��Ǐُ���w�!� ͟��i�)������� +�՟�������ůA� S�e��7���[�m�ѯ y����п+��O�� !υ�7ϩ�����߿�� ϯ�����K���oρ� ��߷�c߉ߛ��Ͽ� #�5�G�����}�=�O� ��[����߲����1� ���g�����f����S��>k�� 3 �k� ����
 ������~��UD1:\&���}�R_GRP� 1?� 	 @��q�m@��������   �&J5nY?�  ���� ���/�//'/ ]/K/�/o/�/�/�/�/�/�/	9�?%?{�SCB 2@�� tq?�?�?�?�?��?�?�?Oq�UTORIAL A���LOv�V_CON?FIG B����	�O[MOUTP�UT C���@���O�O__1_ C_U_g_y_�_�_�_�_ �_�A�O�_oo1oCo Uogoyo�o�o�o�o�o �_�o	-?Qc u������o� ��)�;�M�_�q��� ������ˏݏ��� %�7�I�[�m������ ��ǟٟ����!�3� E�W�i�{�������ï կ�����/�A�S� e�w���������ѿ� ����+�=�O�a�s� �ϗϩϻ������� �'�9�K�]�o߁ߓ� �߷����������#� 5�G�Y�k�}���� ������O�E�O'�9� K�]�o����������� ��������#5GY k}������ �1CUgy �������	/ -/?/Q/c/u/�/�/ �/�/�/�/�/?/)? ;?M?_?q?�?�?�?�? �?�?�?O?%O7OIO [OmOO�O�O�O�O�O �O�O_ O3_E_W_i_ {_�_�_�_�_�_�_�_ o_/oAoSoeowo�o �o�o�o�o�o�oo +=Oas��� ������&9� K�]�o���������ɏ�ۏ���������0�B�,��m�� ������ǟٟ���� !�3�E�W�i������ ��ïկ�����/� A�S�e�w��������� ѿ�����+�=�O� a�sτ��ϩϻ����� ����'�9�K�]�o� �ϓߥ߷��������� �#�5�G�Y�k�}�� ������������� 1�C�U�g�y������ ��������	-? Qcu������ ��);M_ q������� //%/7/I/[/m// ��/�/�/�/�/�/?�!?3?E?W?i?{?�;��$TX_SCRE�EN 1DD��,��}i�pnl/�0gen.htm�?�?�?O�O%O��Pan�el setup)L}�)OjO|O�O�O�O�OXONO�O__ 1_C_U_�Oy_�O�_�_ �_�_�_�_n_�_-o?o Qocouo�o�_,o"o�o �o�o)�oM�o q�����BT ��%�7�I�[�� � �����Ǐُ���t� !���E�W�i�{��������>UALRM_�MSG ?�9��0 ���*��5� (�Y�L�}�p��������ׯʯ����ӕSEoV  �Q��ђECFG Fv�5�1  �%�@�  A��  w Bȍ$
  � �#�5��ƿؿ���π �2�D�V�h�v�]�G�RP 2Gg� 0�&	 ����Ӑ�I_BBL_NO�TE Hg�T?��l�"�0�!s���DEFP�ROݐ%� (%�:ߖ (�a�L߅� pߩߔ��߸�������'��K���FKEYDATA 1I�9���p v��&��ϰ����������,�(�+��$(PO?INT  ]3�5���NCEL_����NDIRECT����� EXT ST�EP��6�TOU�CHU���OR?E INFO OaH�l��� ���9 ]�o ��/f�rh/gui/w�hitehome.pngp��������point�*/</N/`/r/�&  FRH/F�CGTP/wzcancel/�/�/��/�/�/�#�indirec/4?F?X?pj?|?�/� nex#?@�?�?�?�? O$�touchup�?@<ONO`OrO�O$�arwrg�?�O�O �O�O_�8#_5_G_Y_ k_}_�__�_�_�_�_ �_o�_1oCoUogoyo �oo�o�o�o�o�o	 �o?Qcu�� (������� ;�M�_�q�������~ ��ӏ���	��-�4� Q�c�u�������:�ϟ ����)���;�_� q���������H�ݯ� ��%�7�Ư[�m�� ������D�ǿ���� !�3�E�Կi�{ύϟ� ����R�������/� A���S�w߉ߛ߭߿� ��`�����+�=�O� ��s�������\� ����'�9�K�]�������������v��������#5WiC,U�M���� ��<N5rY ������/� &//J/1/n/�/g/�/ �/�/�/���/?"?4? F?X?g�|?�?�?�?�? �?�?w?OO0OBOTO fO�?�O�O�O�O�O�O sO__,_>_P_b_t_ _�_�_�_�_�_�_�_ o(o:oLo^opo�_�o �o�o�o�o�o �o$ 6HZl~�� ����� �2�D� V�h�z������ԏ ���
���.�@�R�d� v��������П��� ���/<�N�`�r��� ������̯ޯ��� &���J�\�n������� 3�ȿڿ����"ϱ� F�X�j�|ώϠϲ�A� ��������0߿�T� f�xߊߜ߮�=����� ����,�>���b�t� �����K������ �(�:���^�p����� ������Y��� $ 6H��l~��� �U�� 2D�V-�X�-�������}���,�/
/�/./ /R/d/K/�/o/�/�/ �/�/�/??�/<?#? `?r?Y?�?}?�?�?�? �?�?O�?8OJO)�nO �O�O�O�O�O��O�O _"_4_F_X_�O|_�_ �_�_�_�_e_�_oo 0oBoTo�_xo�o�o�o �o�o�oso,> Pb�o����� �o��(�:�L�^� p��������ʏ܏� }��$�6�H�Z�l��� ������Ɵ؟�����  �2�D�V�h�z�	��� ��¯ԯ������.� @�R�d�v���_O���� п�����*�<�N� `�rτϖ�%Ϻ����� ���ߣ�8�J�\�n� �ߒ�!߶��������� �"��F�X�j�|�� ��/����������� ��B�T�f�x������� =�������,�� Pbt���9� ��(:�^ p����G��  //$/6/�Z/l/~/��/�/�/�/���+}�������/@?=�/7?I?#6,5O z?-O�?�?�?�?�?�? �?O.OORO9OvO�O oO�O�O�O�O�O_�O *__N_`_G_�_k_�_ �_���_�_oo&o8o G/\ono�o�o�o�o�o Wo�o�o"4F�o j|����S� ���0�B�T��x� ��������ҏa���� �,�>�P�ߏt����� ����Ο��o���(� :�L�^�ퟂ������� ʯܯk� ��$�6�H� Z�l���������ƿؿ �y�� �2�D�V�h� ���Ϟϰ��������� �_�.�@�R�d�v�}� �߬߾��������� *�<�N�`�r���� �����������&�8� J�\�n�����!����� ��������4FX j|����� ��BTfx ��+����/ /�>/P/b/t/�/�/ �/9/�/�/�/??(? �/L?^?p?�?�?�?5? �?�?�? OO$O6O��8K�����aOsO�M]O�O�O�F,�_�O�__�O2_ D_+_h_O_�_�_�_�_ �_�_�_�_oo@oRo 9ovo]o�o�o�o�o�o �o�o*	�N`r ����?���� �&�8��\�n����� ����E�ڏ����"� 4�ÏX�j�|������� ğS������0�B� џf�x���������O� �����,�>�P�߯ t���������ο]�� ��(�:�L�ۿpς� �Ϧϸ�����k� �� $�6�H�Z���~ߐߢ� ������g���� �2� D�V�h�?������ ������
��.�@�R� d�v������������ ����*<N`r ������ �&8J\n� �������"/ 4/F/X/j/|/�//�/ �/�/�/�/?�/0?B? T?f?x?�??�?�?�? �?�?OO�?>OPObO tO�O�O'O�O�O�O�O __�O:_L_^_p_�_h�_�_}��[�}�����_�_�]�_o)of,Zo ~oeo�o�o�o�o�o�o �o2VhO� s�����
�� .�@�'�d�K�����y� ��Џ����'_<� N�`�r�������7�̟ ޟ���&���J�\� n�������3�ȯگ� ���"�4�ïX�j�|� ������A�ֿ���� �0Ͽ�T�f�xϊϜ� ����O�������,� >���b�t߆ߘߪ߼� K�������(�:�L� ��p�������Y� �� ��$�6�H���l� ~���������������  2DV]�z� �����u
 .@Rd���� ���q//*/</ N/`/r//�/�/�/�/ �/�//?&?8?J?\? n?�/�?�?�?�?�?�? �?�?"O4OFOXOjO|O O�O�O�O�O�O�O�O _0_B_T_f_x_�__ �_�_�_�_�_o�_,o >oPoboto�oo�o�o@�o�o�o��{��������ASe}=��sv, ���}����$�� H�/�l�~�e�����Ə ؏����� �2��V� =�z�a�������ԟ�� ��
���.�@�R�d�v� ���o����Я���� ���<�N�`�r����� %���̿޿��ϣ� 8�J�\�nπϒϤ�3� ���������"߱�F� X�j�|ߎߠ�/����� ������0��T�f� x����=������� ��,���P�b�t��� ������K����� (:��^p��� �G�� $6 H�l~���� ���/ /2/D/V/ �z/�/�/�/�/�/c/ �/
??.?@?R?�/v? �?�?�?�?�?�?q?O O*O<ONO`O�?�O�O �O�O�O�OmO__&_ 8_J_\_n_�O�_�_�_ �_�_�_{_o"o4oFo Xojo�_�o�o�o�o�o �o�o�o0BTf x������ ��,�>�P�b�t����]���]�����ÏՍ����	��,��:��^�E� ����{�����ܟ�՟ ���6�H�/�l�S��� ����Ư���ѯ� � �D�+�h�z�Y���� ¿Կ�����.�@� R�d�vψ�ϬϾ��� ����ߕ�*�<�N�`� r߄�ߨߺ������� ���8�J�\�n�� ��!����������� ��4�F�X�j�|����� /����������� BTfx��+� ���,�P bt���9�� �//(/�L/^/p/ �/�/�/�/���/�/ ? ?$?6?=/Z?l?~?�? �?�?�?U?�?�?O O 2ODO�?hOzO�O�O�O �OQO�O�O
__._@_ R_�Ov_�_�_�_�_�_ __�_oo*o<oNo�_ ro�o�o�o�o�o�omo &8J\�o� �����i�� "�4�F�X�j������ ��ď֏�w���0� B�T�f������������ҟ���� ���>� ���!�3� E��g�y�S�,e��� ]�ί�����(�� L�^�E���i������� ܿÿ ����6��Z� A�~ϐ�wϴϛ����� �/� �2�D�V�h�w� �ߞ߰��������߇� �.�@�R�d�v��� �����������*� <�N�`�r�������� ��������&8J \n����� ���4FXj |������ /�0/B/T/f/x/�/ �/+/�/�/�/�/?? �/>?P?b?t?�?�?'? �?�?�?�?OO(O�� LO^OpO�O�O�O�?�O �O�O __$_6_�OZ_ l_~_�_�_�_C_�_�_ �_o o2o�_Vohozo �o�o�o�oQo�o�o
 .@�odv�� ��M����*� <�N��r��������� ̏[�����&�8�J� ُn���������ȟڟ i����"�4�F�X�� |�������į֯e������0�B�T�f��$�UI_INUSE�R  ������� � g�k�_MENHIST 1J���  �( ����*/�SOFTPART�/GENLINK�?current�=editpag�e,ZAD15,A1���-�?��(���menu��153ϛϭϿ����߿��1��!�3�E�W������2ߥ߷��� ��j�|��(�:�L�^������4���L����'t�v�2�-�?�Q�c�^����48,2h������������۱��
.@Rdv �� �����+= Oas���� ��/�'/9/K/]/ o/�//�/�/�/�/�/ �/�/#?5?G?Y?k?}? �??�?�?�?�?�?O ��1OCOUOgOyO�O�O �?�O�O�O�O	__�O ?_Q_c_u_�_�_(_�_ �_�_�_oo)o�_Mo _oqo�o�o�o6o�o�o �o%�oI[m ���D��� �!�3�O<�i�{��� ����Ï������ /�A�Џe�w������� ��N�П����+�=� O�ޟs���������ͯ \����'�9�K�گ \���������ɿۿj� ���#�5�G�Y�D�� �ϡϳ��������� �1�C�U�g��ϋߝ� ���������߆��-� ?�Q�c�u����� ��������)�;�M� _�q������������ ����%7I[m�j��$UI_P�ANEDATA �1L�����  	��}/frh/g�ui�dev0.�stm ?_wi�dth=0&_h�eight=10�� � ice=TP�&_lines=�15&_colu�mns=4� fo�nt=24&_p�age=whol�e� �h�)prsim/X  }[������ ) ���#/
/G/Y/@/ }/d/�/�/�/�/�/�/�?�/1?h����     ][�in?�?�? �?�?�??�?_O"O 4OFOXOjO�?�O�O�O �O�O�O�O�O__B_ T_;_x___�_�_�_�_E7 � �U�Oo$o 6oHoZolo�_�oO�o �o�o�o�ouo2D +hO����� ��
���@�'�d� v��_�_����Џ�� �Y�*��oN�`�r��� ������!�ޟş�� &�8��\�C�����y� ����گ�ӯ����� F�X�j�|������Ŀ ֿI�����0�B�T� ��x�_ϜϮϕ��Ϲ� �����,��P�b�I� ��mߪ��/����� �(�:�L��p�㿔� ���������U��$� �H�/�l�~�e����� ���������� D V���ߌ���� �9
}�.@Rd v������ //�</#/`/r/Y/ �/}/�/�/�/�/cu &?8?J?\?n?�?�/�? �?)�?�?�?O"O4O �?XO?O|O�OuO�O�O �O�O�O_�O0_B_)_`f_M_�_�/?}��_@�_�_�_
oo.o)�_ So�5Boo�o�o�o�o �o@o�o�o!W >{b���������/��83;��$UI_POST�YPE  5�� 	 �;���a�QUICK�MEN  p�����c�RESTO�RE 1M5�  ��*defaul�t�;SING�LEԍPRI�Mԏmmenu�page,148,2 1<�q����� ��J���П����� ��<�N�`�r����"� �����ϯ��
��.� @��d�v�������O� п�����ï%�7� Iϻ��ϖϨϺ���o� ����&�8�J���n� �ߒߤ߶�a������� Y�"�4�F�X�j��� �������y����� 0�B�����a�s���� ����������,> Pbt��������SCRE��?���u1s]c�u2!3!U4!5!6!7!�8!�TATl��� ă5Y�USE1Rks#�U3�4�5�6��7�8�a�NDO_CFG Np���P�Qa�OP_CRM5  �U&a��PDd���None���_INFO 1O55f 0%��/ �8o/�/�/�/�/�/
? ?�/@?#?d?v?Y?�?�?�?�?��S!OFF?SET Rp�j!�?����!O3OEO WO�O{O�O�O�O�OO �O___J_A_S_�_ w_�_�_�Kŏ�]�_
o�
�_/o�8UFRA�M%�/P!RTOL_ABRTSoN#kb�ENBtoehGRP� 1S����Cz  A��c�a��o �o�o�o"v,>�cj��U�h#!�kMS�K  �ef!�kN6Pa%^)�%�_���e_EVNs`�t�&�v�2T�;
 }h#!UEVs`�!td:\ev�ent_user\�7�C7<�o� YFq�/�SP5�:��spotweldl�!C6��r���#�t!�K�	�>�� q��-��q���Q�c� ܟ�� �����ϟH�� l��)�_�����د�� ��˯ ��D���z� %�����[�m�濑�
����Ǻ�WRK 2U�a8�nπ� \ϥϷϒ������� �#���G�Y�4�}ߏ� j߳��ߠ���������1��B�g�y��$V�ARS_CONFuI�V�; FP�����CMR�b2�\�;xy� 	�$ ��01: S�C130EF2 Q*�	����X�ȸ�p�  #!?��p@pp"p�z� o]�g����@����������`�u�A����,�? B���G� K��l���_�� �����2� hSe�Q�����IA_WOF�]<^-˶,		�Q;%|/+'G�P �> ����RTWINU_RL ?�������/�/�/�/�/��/�SIONTM;OU� ��%��^S۳�S���@�a FR�:\�#\DATA�؏  �� wUD166LOGC?7  \9EXh?'q�' B@ ���2{1U��?{1�?��?θ � n?6  ������2�zt�`F��  =���BA��?@>|=TRAIN�?A4QB�d�CpBEFF�/B�0�(��_� (��I�M��O�O�O __P_>_t_b_|_�_��_�_�_�_�(_GE23`�/C�
�`'pX4b
g�0RE!0a�i\���LEXdb�����1-e�/VMPHASE  ����C ��RTD_�FILTER 2]c� �&��T� �o+=Oas �����o�������1�C�U�g��)S�HIFTMENU� 1d�K
 <b�<%�?ŏ2���� ɏ�ُ�8��!�n� E�W�}��������ß�՟"���	LIV�E/SNA��%?vsfliv�n4����# SETyU��W�menum��r��ѯ�"��3e�`+|�MO3ftn�-z��ZD�gQm˳�<�A�P�$WA�ITDINEND�8L!�k�OK  !�醼 :��S����wTIM5���Gr�͔�%˴��ӿx�򿆸RELE�a�5��k��/6m�_ACCTJ�4� !��_?17 h��%�5�<����RDIS��ο�$XVRna�itn�$ZABCv��1jQk ,�@r�2=��-ZIP2kQo���)����MPCF_G 1l��l!0L"��q�7�MP��m����P�������`�~*�  6n�G��6�"IG�o�5�j�5�i���A�H�C�/��CQ�Ch�<�0�Q���;�=�/";��P������ɿNO?��������������6�?6W�lT����5@�?���,�����p9�������C��C�0B������G�Ҫ�9lw7³���,I�䮵9lfw$@�PJ \r��������A6�����J�p`n���_CYLIND��aoR� �p6? ,(  *o��w3l����  ��//'.iJ/�n/ U/g/�/��/�/�/// ?�/�/F?-?j?Q?�/��?�?�Cp*� �g��?L^���6O@!OZO?I�?�O?G��A�A�=SPHER/E 2qO�?�O T?�O_�O:_�?�Op_ �_�/�_E_+_�_�_ o �_Y_6oHo�_�_~o�_ �o�o�o�oo�o 6��ZZ�� ��