��   2�A��*SYST�EM*��V9.1�0185 12�/11/2019� A 
  ����PASSN�AME_T  � 0 $+ �$'WORD�  ? LEVEL  $TI- 7OUTT��&F�/� $S�ETUPJPRO�GRAMJINS�TALLJY � $CURR_�O�USER�N�UM�STSTO�P_TPCHG �V LOG_P NeT�N�  6 �COUNT_DO�WN�$ENB_PCMPWD� �$DV_� I�N� $C� CkRE��A RM9z� T9DIAG9�(�LVCHK| FULLM/�YXT�CNTyD�MENU��AUTO+�FG�_DSP�RLS��U�BURYB�AN�!eENC�/  C�RYPTE �� ���$$CL�(   ���TK!��	��	@ V� �IONH(�  �i\!IR�TUA� J/�$D�CS_COD?����O%�  W�'_� �/�(S  J�*�� � �&�A�91�"�!	 $R!�� =,? B?P?f?t?�?�?�?�? �?�?�?OO(O>OLO�bO��3SUP� �:�dOvO3F�O�O�O��  !\Q��&_ ��� V�[t&W��j��T�O ~_��<W:_��t �V�U��Y�ELUGH 1}�) t �)oo'o9oKo]o oo�o�o�o�o�o�o�' �_	-?Qcu �������o� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ ������/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ������� �� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ������
��1�C�U� g�y������������� ��	�-?Qcu ������� �%