��   :�A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����FSAC_�LST_T  � 8 $CLN�T_NAME �!$IP_AD�DRESSB $�ACCN _LVL�  $APP~P  ���$8 �AO  ����z����o VE�RSIONw  �i�?IRTUALw�'DEF\ � � ��� ���ENOABLE� �������LIST 1� �  @�!�,��)��� (yL^���� ���-/ /Q/$/u/ H/Z/�/~/�/�/�/�/ �/?�/:? ?q?D?V? h?�?�?�?�?�?O�? 7O
OOmO@O�OdO�O �O�O�O�O_�O3__ _U_<_z_`_�_�_�_ �_�_�_�W