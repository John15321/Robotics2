��   T�A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ������DMR_�SHFERR_T�   $�OFFSET �  	��/G�RP:� �$MA��R_DO�NE  $OT_MINUSJ 7 	sPLzd�COUNJ$REYFj�PO{���I$BCKLS�H_SIG�E?ACHMSTj��SPC�
�MOV�n ~ADAPT_�INERJ F�RICCOL_�P,MGRAV8�� HISI�DSPk�HIFkT_7 O ��Nm�MCH� S��ARM_PAR�AO dcAN�Go y2�CL�DE7�CALI�BDn$GE�AR�2� RINYG��<$]_dΗREL3� �1  	��CL|o: � ��AX{  $PS�_�TI���T_IME �J� �_CMD��"FB�VA �&CL_OyV�� FRMZ�$�DEDX�$NA� %�CUR�L�W���T{CK�%�FMSV��M_LIF	��'83:c$�-9_09:_��=��%3d6W� �"�PCgCOM��FB� yM�0�MAL_�#ECI�P:!o"7DTYkR_|"�5�:#�1END�4���o1 l5M̦P PL� W ݀�STA:#TRGQ_M��� KNiFS� uHYsJ� hG�I�JI�JI�D���$�ASS> �S���A�����@�VERSI� �G�  �i~�AIRTUAL�O��AS 1�H� ��� 	 ��\_G_�_k_�_ �_�_�_�_�_�VP���em�U�ABo0l���'R��� ������X����2�/o�ooUl��o�o�o�o�o�k ;Ar*gyd����d������=L3����?����@�=�b�t������� ��Ώ�����(�{ US�a�K����D  2���ğ֟蟀����0�B�T���< ��~�������Ưد� ��� �2�D���Pr�(�x���������� �Ͽ���>�)�b�`Mφ�qϖϼ��$4� 12\���N���MlD�L����E�� O���M�9:���@�|vA��|�@�-�32��:�;�;�����B�  @ߙϽ��y�dߝ߈�A��:�߯���߈�� ��9�$�]�o��LLêK��X���� ���T���P�������'���%��345678901G�O�t� x�q���m��������� ��D�}���z�H ��lZ|����� .��2 Vh ����n@�� �/r�U/���/ /�/�/�/�/8/	?? n/�/N?<?r?`?�?�? �/�?"?4?�?�?O8O &O\O�?�?�O�?�?�O FO�O�O�O"_xOI_[_ �O_�_|_�_�_�_�_ >_ob_t_�_�_Boxo fo�o�_o�o(o:o �o,<b�o�� �oP�����(� ~O���.� ����� ��܏2�D��h�z�H� Əl�Z�|�����ɟ۟ .������2� �V�h� �������n�@�¯�� ��r���U������� ��������8�	�� n�пN�<�r�`ϖϨ� ����"�4Ϯπ��8� &�\�n�}��ϕ�����,[�����9��$�PLCL_GRP� 1S��� D�?�  ���;��_�J� ��n��������� ��%��