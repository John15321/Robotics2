��  	w^�A��*SYST�EM*��V9.1�0185 12�/11/2019� A  �����AAVM_�WRK_T  �� $EXP�OSURE  �$CAMCLB�DAT@ $PS_TRGVT��$X aH]ZgDISfWg�PgRgLENS_CENT_X��YgyORf  � $CMP_G�C_�UTNUM�APRE_MASwT_C� 	��GRV_M{$�NEW��	ST�AT_RUNAR�ES_ER�VTSCP6� aTCb32:dXSM�p&&�#END!�ORGBK!SMp��3!UPD�O�ABS; � P/ �  $P�ARA�  ����AIO_wCNV� l� �RAC�LO�M�OD_TYP@F+IR�HAL�>#�IN_OU�FA�C� gINTER�CEPfBI�I�Z@!LRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CESI0�!H1�!"PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W� @V�R!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2 � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1 UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t�cbMO� �sE 	� [M�s��2�wREV�BILF�?  �AXI� %��R  � O�D}`j�$N5O`M�!b�x�/�"u�� ������`��@Dd� p E RD_�Eb��$FSS�B�&W`KBD_S�E2uAG� G�2B "_��B�� V�t�:5`ׁQC �a_E�Du � � �C2��`S�p�4%y$l �t$OP�@rQB�qy�_OK���0, P_C� y��dxh�U �`LACI�!��a���� FqCOsMM� �0$D���ϑ�@�pX��ORB�I�GALLOW�� (KD2�2�@V�AR5�d!�AB ��BqL[@S � ,K�JqM�H`S�pZ@M_�O]z���CFnd X�0GR@���M�NFLIx���;@UIRE�x84�"� SWIT=$�/0_No`S�"CFu_�G� �0WARNMxp�d��%`LI�V`NST�� COR-rF�LTR�TRAT� T�`� $AC�CqS�� X�r$�ORI�.&ӧRTβ`_SFg CHUGV0I�p�T��PA�I��T�!�|�� � �#8@a���HDR�B���2�BJ; �C��3��4�5�6�7b�8� � ����x@�2 @� TRQ��$%f��ր�Ǎ��_U����e`C=Oc <� ��දȨ3�2��LLE�CM�-�MULT�IV4�"$��A
2FSN�ILDD�
1R���z@T_1b  4� STY2�b4�=@�)24����E��� |9$��.p���6�I`�* \�T�O��E��EXT����ї��B�ў22��0D��@`��1b.'�B ��G�Q� �"Q�/%�a���X�%�?sdaD�U�  Sҟ�;A�Ɨ�M�� �� CՋO�! L�0a�� X׻p=Aβ$JOBB����ֈ�TRIGO�" dӀ�����X�-' x���G�ҧ��C�`�.�b# tӀF� �C3NG�AiBA� ϑ ��!���/1��À�0����R0P/p����$
�|��BqF4]�
2J]�_RN��EC`J`�e�J?�D/5C�	�ӧ��@ʤ�P�O3л!% \�0RO�6� ��IT�s� NOM_ 8pn#�c ���kTU�@P� � ���&+P��� ӨP�	ݭ��RAx@n �3x�A���
$TF3�%#D3
T��wpU(�13�}�%mHrzT1�E���ޣ��#ݤ�%ߢQlYN�T�"� DBGDEf�!'D�]�PU��`�@t����"��AX���"�uTAI2sBU�Fۆ�0>"�1( ���P&V`PI84'*mP�'M�(M�)B ��&F�'SIMQS��@ZKEE3PAT�zЙ8"�"<!_MC��)S�0��`�JB���ľaDEC�g:� g5���* ��U�CHNS_EMPͲ$G��7��_��c;�1_FP,)�TC�6S���5@�`%��4�} ��V�����W��JR����S_EGFRAq�O��| #PT_LIN�KCPVF�� �C$+���ckBZ�PBzr�g��@6,` + �Ԧ��A�0��Ad0�o`Ar�D���Id1SI!Zh���	T�FT�C�Z1Y�ARSm��C P@'�Ic\1@cX�0<@�L����0�VCRCߥ�sCC���U1@�X�1��2�Mpq�U�1`�X�Q�UDݤأiCk�p*�
DK`݀fL��RhEVRf �Fha_	EF�0N�f�Pd1�&h��5�jC}�=+�VSCA[��IA�fgC13��-�y	�ׇMARG��D�a�F@@���1DcQ��r�0LEW�h�@�R�P<��o�l��RɄ.� ����ǯ��� 5ڡR�`HANC��$LG5��a�� Ӑ��ـF��Ae����0RYr�3
�����
�@ �RA��
�A�Z�0Q�N`�O��F#CT��sp�F��R��0P0b ADI��O ��+���+���&���5�5����S[�g���'BMPUD(PY�1���AESCPjc��W*��N  SuU0ۑuU�/)�TIT'q�<�b�%ECA:!�!E'RRLd��0�&Q��OR�B$������~��$RUN_O��SYS��4������u�REV�c��?DBPXWO�P�=1d�$SKo�"��DBT�pTRLn�2 �C AC��0��%�m�U DJ�p��_p�!A�ǀM�P5L�A_2WA��j�EE��D!w�!%R|hO�UMMY9��ڠ�1� / DBd[��3���!PR�Q� 
�ٱ9��4� г$α�$ Q�Lة5L�z����6�^zd�PC�7*�~ze�PENEC0�Tq8I����R�ECOR$�9H� m��4$L��5$أ�"E���R@���VA��_Dց� R3OS �"SK������I�=�א��PA���JVBETURN,���SMR(�U #�CRʰEWMDB�0GNALV �"$�LA� [�*6$=P-�7$Pv�s�#8o�!�PC��#�DO^@-�Ŵ���R>˶GO_AW�ܱ�MOz��p�O�C_SS_CN4�YO��:��T��0���IDT�T�2��2�N���O@�J��v`Iְ ; P $>�RB�B��PI�P=Ol�I_BY��v���TVR��HNDG$�< H�`�1a�x@cS��DSBLI���s���0}���LS�$�=��0� ��FB�FEձL�9�����5��>D�$D1O�1�C�pMC�0q��4��9�RH��W8��K4ELE�urz�C��SLAVr?xBINS ���#��:��_R@P�@\` �pS�}�l�}�l�{u��D[!e��ے�I�Ȋ�B��W��D�NT�V�#�VE�$��S�KIlA4;3��2�UB�1J�f�1C�
DS�AF7�5��_SV>6�EXCLU-���XrONL�0Y�Y��s����HI_V�Հ�RPPLYo�RbCsH� �0_M�}Q�VRFY_I�z.Mms$IOv0���}��1UB���O�j�3LS����4�!��:@�P��$�ĆAUTOCNE ����.�N�GCHD�s��_��l�3s�AF��CPe�T!��р� #Ao���_�0 w ��NOCtIBxB�pT��A ܢ��_SG�` �C � 
$CUR8�U��!" �� ��B�����ANNUNC�#������b���()%!��-*�I&�EF��IC�D� @�F
"a��POTX�aө�������j�� e M��NIߢ!E�·"�G� A��$�DAY��LOAD�`Ԟ��"��5����EFF_AXI�%Fo�%Q�O0���:�_RTRQV1GC D�a��?0�RK3x�0S45 2Fz@8]w:1a��A0p/1NsAH 0B!�1A�T��2�ûvDUX��u�.�CABsAIs"�p�NS�1�PID�@P�WSs�5�AWpV`�V�_�0q0�P�DIA�GysAJ� 1$VX��ET	`�UrT��EJ��{RRf��!�T�VE�� SW�|AZ�sP�0�:5q0G�}P:1OHP5�1PPL|@�SIR|�{RB�P �2�3%qZQC �BB���H�^��E`��5q0I�$0?0���URQDW&�EMSB�?UA�p�E<jB�TLIFEpK#iP��uRN|QFB�U%!�zSFB�a�%"C����N��Y'p�F3LA�t& OVڰ�V�HE��BSUPPIO(��uRI�_�T��Q_X�d�� gZjWj� g��%!���6�XZ*�ϡfAY2xhC��T��DEQN�pBE%!J�� �F�_8p�A���p�K{ `Q�CACH�*r�bSIZ�V�Pz`�N��UFFI`�oP�ў�2���6���M;��tL �81 KEYIMAG �TM��!�^q:��Yv����OCVI9E�@�qM $0���L~��;�?� 	���р�dNG0��ST��!�r���t����t0�t0�pEMA�ILo����!��5FAUL�"O�r��/�N��COU���T��~)AP< $9��p�S�0�0IT��BUF�g;��gE�o�e�%�PBe�p�C:���8:�|�G�SAV��r��[@�b��@ˇÐ)&P ��p印�D��_e����� �OT겮�3P`m ��0�z3�AX���f x Xe�C�_G:|S
� YN_�A��Q <�Dk�O���U�BM�2�PT� �F�$�DIB[E7�����R��$ G���!&�Ǳ����c :�9�S�0���-��C_ᰤ�AK�$�����RVq8���DSPnv�PCe�IM��\���<�3@U9��P�] �IP���A�`[�CTH�`3�O�0T��\�HSȓ>�BSC���`e�V��
�\�X���*4NV��G;����`Y�e�F|A}�d0>���Z��SC%Ba���MER)�FBgCMP)�ET�� TLrFU`D�UY���R�mb�CD�R�ܠ'�"�e��N)O�n!UG0*���H�%���%P���C�
ō-"�!��:��o VH *
�L ��)�9���G ��� }�Z{ƥ!{�1{�1�{�6q{�7x�8x�9Px�|PzȄ�1��1��U1��1��1��1��U1��1��2��2�˪��2��2��2��2���2��2��2��3J��3��3�˞�3��U3��3��3��3��e3��4��2XT6An!W��߸���V��u�蟐����`FDR^%DXTE�V� �.�uR�
�uRREMr^@F���BOVM5�z*�A3�TROV3��DT��S�MXb�I�N3��PR�"AIND�q�cB
��ɐ}���G@e��C\�p�UkADO6�\�RIVW�R�BG�EAR5�IObEK#�cDN��1`X� �zp`dCZ_MCM�p`uQ �F�PURζ�Y ,���?3 �P>?o {A?oE� w���������Z� *PPM�2@RI��0r��ETUP2_ 3[ 0q�TDʠ�1p�T�����qr�wBAC��\ T�pr��)�%w#@ó�TIFI�A����d���@/PT�B�FL{UI�t] �@�x;�UR�A���R��Б
��:C_0I�$��S_?x�J��CO��"�VRT|��� x$SHO^14 #�ASS�-��U̠��BG_ �!.��!��!��!��FO�RC�hDATAZ)A^�rFUZ1���]#2���j�`)A_� |��NAV=�S�����S�~�S$VISI��6��SC=�SE� ���5V� O�1&1B�F�4@�&$PO�� I�A�FM�R2��`  ���2���6�@!3J�)�CE#�_��9��_@IT_Yִ�]@M������DGC{LF�EDGDY�8LD���5�V���TR�M���sa��v9? T�FS
��t�b P��RB��}��$EX_RAiHRA1PY�X��RS@3�K5�Fs�G&�	5c �� ֳ�SW��O0VDE�BUG$�A(�GRt� opUz�BKU���O1M� �0P�OZ0Y�@���E�@M��LOOM�9QSM0E��J���P_E� d rp��T�ERM[UedUua�l�ORI֑`Pf~dV�SM_㐄�`PgdU��Q �Xh�dV� UP�ri�3 -���2d�rS��Pe� G�Z @EL�TO���A�FIG�bZ �Agp�T�T�f$UFR��$��aM`ѵ�0OT�ZgA�TA��lcN;STאPAT��`��bPTHJ�ϰEp�p�ذbART؀�"e)�؁���REL<�j�SHFTӢ�a�h_�R��̳�V% �P$�Wph�1�8���t�SHI�`�4�U � ҁAYLO ��m���l� ��a}!�ޠERV��Sq� x��hgא�b �K�u�.�KRC��AScYM���WJ+g���E��a�y�ұU�א���e@�v�eaP��ppE�2vORא�M3fGRJQ
4j�X"�B0V�`G`l�� H9O�6Dk ��aN,� �OCaQ@$OP�$e�i�F�����2ՀRY��aOU��c�PTR�e����a��e$PWR��IM��rR_˃�d� ��P�cUD��cS�Vl���֔l� $�H�!��ADDR
��HMQG�b����������R�"1m H��S���! ��.����畫�SEz1�#��ySܰ
3n $Z �À_D��P�.�P�RM_�"����HTTP_��H�1o (��OBJ�� ��)$��LE�yc��d�p � ��睱AB_��T�@S��S���{KR�LK�HITCOU � À�!퀶���0��M�SS��v��JQUERY_F�LA!a��B_WE�BSOC�"�HW���a1q�7�IONCPU�B�!Ou� ˡ�Č���������¿�IOLNr� 8��R	� $�SL2$INP7UT_PQ$�ܸ�P�# ��SL]A�1 sðٿ����s��rNAIO^C�F_AS8Bt�$L&��&q �!]�/a�ɳ�@ҳUp�HY���lïAG�U;OP5Eu `X�������ā������P �����������UQr� M�qqv lq@�;sTAkr��A�T�I��.�a�Z0S��`PmSR�BUZ0ID~0 ��z���y�lQ!�u�&z`w�3�f�G���N��Z0���IR�CA��� x �Ĩ��CY�EA{���!���%�¦R�`�q|�8�DA�Y_��}�NTVA����i�¦eu�i�S3CAepi�CL���"����� qy����X�b����N_ՀCQ�Ђ�W�rz�O � �������y�G�]�O!� 2y�)q{pP���P�LABza�n�Z0t�UNISb�PITY��"ѳ�&�IR$6D|�R_URL� �$AL10EN�@�� t�PH�T�T_U�� �Jt�q} X ��t�R��" "�0A�D�,J�8#FLt@�80
K�3�
�UJR	5~ ���F|@1w�Fgw�D��$J72�O^!�$J8�	7�@H\��7s�� 8�	ޡAPHI@Q���Df@J7J8��
L_KE�� � �K��LM���  <��X�RK��� �WATCH_VA�!pp��_FIELD��y`�L&��� �0paVyp�ֆCT��E��B�R�LG����� !��LG_SIZ���@�3@�,O��FD�I�� ,Q��]P���� J&3@J&O�J&�J&]P�J&�q�E`1_CM ^c�!{@�*h1F��'��$��(�#r��&3@�&O��&��'I�(�(,P�&]P�&��RSI�`  M(�PLN��B�����@{A�g1���K�u1��L~3t2DAU�5EAS������2Ʀ0GH���Q[�BO�Oܑ�� Cr�[�IT8��4<`n�sRE(��8SCR� ,ڣs�DIm�SG`G@7RGIPR$D/L� f�քYB��[�S��Z��W7D[��4f�JGM��GMNCHH�[�F�N�FK�G��IUqF�H2p�HFWD�H�HL�ISTP�JV`�H�P�H�0�HRS3YHJ��Kc�C4tS�f�x�kG�YUJ��DjG  3yE�{��BG�I�`PO�WZ&ES�"�D�OC���FEXb�TUI�EI/ ���/! �dDa�CNc�@��p��� 4	��EpANO�GfANA[�ā�A�It瑜��DCS�Z���c���bO�hO"�gS?��b�hS�hNHIGN�����A��(��dDE��pTLL �q��|A��*Є���T�"$���}��Դ��SA����@��ʰ��Z�� �P1�u2�u3�qL��R�`*�G� ���V��c� �5�z�x�6��P�6�V.�ST��R�0Yy���`Q� �$E_�C_�� I�n������T)ч Lo�������x������_�EN�S�_���pBC_ �L���X���@���MCh2� =���CLDP��TRQLI��D�2�FLGZ�2�3�f�b��Duf�`�LDf�P�f�ORGjQy�~�(RESERV���Ŕ��Ŕ� #�3�� � 	O�jUA�Ff�SVX0D�R	����'�RCLMC�5�şןG���'���M�ՠJ�/�3$DEBUGMAS�ÐS�D�"��T�`p�Er� TZ��FRQ���� � �H_RS_RU�ځ��A)��UFREQ�� J�$``�OV�ERh����v|Pn�AEFI��%�������ӡ� \8 ��$U��g?����PS�p
7 	�C�06�BҒ��G�U�Н�?( �	bMISCi�� dq1�RQ5	f	TBB@�� ��aa�AX9�!	�"�EXCES��P۳)M��.����9��"ܲSC� � H���_G���,�P�� �2��K���|�أB@��B_�FL�IC��B@QUI[RExSMO��O���d�"�L܀M��� �
��19Э��5��`pMND�1e�/��o2f2�x�D�#�4I�NAUT(A�4RSM� ��pNZ�b!�Sx^�pe�PSTL.w� 4��LOC��RI1P�EX��AsNG�b�� T�b -Aե��p�x MF�%7�+�ۂ�|@�e�c0��SUP~����FX/ �IGG�1 � ���ۃb!Cۃ�Vۄ ��V�P���R���R���`���SD�w��TIjȻpM�b!M ��� Mt-�MD*��)8��`C�L�@�H�C�GDIA�D�2 W]APC��q��C�D�3)���MOh�/� a�CU�V�����$�PA_��.� �`/��7㉠f��
 B��P��>P���P���KE�RR�#-$B8�����ND2N�N�D2_TX�XT�RA�cp`��9�L�O�0/�_��	�i2�����q�MRR2൜�� -��1A$� ?d$CALI��c%�G�a�2�pRIN��!�<$R� SWq0S� `�ABC>�D_JV ����7�_�J3K
E1SPH���PEl3k(�񱀦��J`��4��OiqIM`�ŲCSKPS��� �c�J�1ŲQ�%�8%'�_AZ#���=!ELNq�N�OC�MP�Ʊ��z0RT��h#�1�����1��(o`�*Z�$ScMGMP�n�JG��SCLB���SPH�_�`Ű+0�#\ ���� RTER���`� _�`�*�A0P@G�Ų4DIS!�"�23U�DF�pv<1LWB8VELD��IN�Z`e0_BL �`��m4���J]4r7�7�4ϠIN� ���!���5QB��
�1��_̰ ��5�2#5�N��4z�936p�D�HB�r ����p$aV� ���#oa$� X����$\���R�����H ��$BELN ��!_oACCEs1 �H<`��@IRC_0����NT��/�$SPSB�7�L�p� �DL��0�G3�`�F;�I�G�C�G3�B��E�_�qPB-P3Q����A7_MG��DDPQ2��FW����ClU�C�BaXDE�[PPA�BN�GRO� EE CR�q�_D�!�q������A�p$USE_t� �cP�CTR�d�Y�Pb@"� ��YN�߰Aa`f�Z�aM����bJPO_0�AGdINC���RpT¸ig��ENC0L���A�B��@IN�7�I�B�e��$NT|]3�5NT23_@2���cLOQ0���`-�IP����fF0����� ����e��C�0�fMOSIUQ����3Q�ŲPERCH  s+�2 ]w�hs��r n���c'["e
P2P�	A'R�uL�T������e��z�vvTRK�%ʁAY��s��,� 'R;�0��n&��wbȠMOM��»������S�G��C�R� �DU�(RS_BC?KLSH_C'R�� ��<v,�"c��݃�b�|1a%CLALM�dp��m�@�CHK�|�NGLRTY�� 5�d����_Z�1t'_UM��l�C��^Q��!����LMTh_AL��V#��j�E�� Ð�����E���H}����r��xPCnq�xHp���TUl�CMCv\^PbWCN_�NuLc��SFtA�yVb��g�!8�'R��<�CATs�SHZ��bT �f]����f��A�	� fQPPAs�gb_Pr�V�_�� 3�Qp�C�U�F�JG>�X�I�K0�OGV�2TORQU�P�/sL��P��Gr1�P��_W��,��!@QAٴBCصHCصI�I�IHCF$�˱�X-��ZPVC�@0����N�1T�RPh�$!ZƇJRKT̙ƴ�D�B� M���M��_sDLBA�rGRVߴ`��BC��HC��H_�8���@�COS�p �LN��6�W�=�B@ 8ٵ 8�
�t�b�(���1Z1�Gv��MY?Ѳ���='���THET=0uNK23HC��l<C@�CB�CB<CC� AS�'�
�5�BC5��SBBCS��'GTS��QCo/���'��'��q�$DUC��w���t5��5eQ�q_��NE��AKS�z)!8 @�сA���'����LCPH����e��SW� o�b�o�q���֙�����V@�V5�2@X�UVg�Vt�V��V��UV��V��V��H@�@Y�_W�ܡvt�H��UH��H��H��H���O1�O@�O�	V�O�g�Ot�O��O��O*��O��O��F��"��~bՃ3�SPBA?LANCE_�Ѯ�LEj�H_��SP��1S��b��q�PFULC�"�"q���:1�|!UTO_<>�F�T1T2B)�B2N%��B�`b$�!f�� ���B}C��T�pO�50�AɰINSEG�B qREV�& p�agDIF��91��'6321�	�OB�!	���Ó�2���`0���L�CHWAR�R7BA�B%���$MEC�H+���9a?1T�AX�9�P�X6�#B7 �� 
Y2��{A�eRO�BQpCR'R�5M�� �CyA_A�T� � x $�WEIGH6`��$1��3X�I6a�`I9F�QjPLAG'b�qS'b� 'bBILEcODo�#p�2ST�@"�2P�!	��0`@Ơ�1�0��0
�`yB(a�A�  2�.t�6D�EBU�3L�@<B���MMY9�E� N8��D�$D�Axq�$�@S��� ��DO_�@A�1� <�0VFL U�$(a�B&B@N�c�H�_p(`CBO� ��� %��T��`�a��T�!~D�@TgICK�30T1�@%NS��WPNQp1 �CQpRԀ(a!2iU!2uU��@PROMP6cE~� $IR���&aL��R�p�RMAIо�aa8b�U_@��S� B�:`R��CO�D[CFU.`�6ID�_ppe� �R�G_�SUFF
� hCa�QdRDOlW0� mU @lVGRC!2 Id�SUd!2`e!2le���Id�De@��0H� _�FIZA9�cOR�D&A �0�B36���b&a�@$ZD�Te\�CA�E�4{ *�!L_NAQ�WPriUDEF_I )xr�V5tuU-BhV7D`hVasuUou�VIS��@���A��hT�suS3tD���D4l���7BD5 (���t[CD��O��BLOCKE�Cci_`{_�W�qIbC`UMHe rIdasIdouId�rUb K�TeDsUdtUb5F�� �q`c,0B�`er`eas `c���EhPP� �t,P�q��@W*�)� ����TE���D� ALOOMB_C�^�0�2wVIS!�ITY�2�AS�O'CA_FR1I2#��� SI�q��B�RTP��_P��3tC
�2W��W��������9_��jaEAS�3jb@d������p�R��4���5��6�3ORMU�LA_I��G�	w� h �N7��ECOEFF_O ;Q� ��;Qr�G��3S�0�BCA �O�C�CAGR�� � �� $ �u"�BX+PTM�� �AR(�,%��CER� T	�tne@�  +"LLkd:�pS�_SV�tw�$L�e@���v�e@�� ��SETU�sMEA�P(`F��0�CA�b�0� � ���0 �@o��Q2��q�rWP�q�	�tբܑubÕQ��p�q�p+���� ��PREC�a�0��MSK_���� P�11_USER^!�"}�0��}�^!VEL"�}�0��r!1I�`J �MTQ�CFGs��  �YP� OG2NOR�E�0P���0��� 4 ݳB7�2H1XYZ�cJ!o yCzH0 ��_ERR�1C� �I�Q�Pۣ�@�aAi����@BUFINDX�po wMOR� H�0CU@�QH1���Q�ax���"�a${0���~q�E@;���G�� � $S�Ij����P�!��VOx����0OBJE���ADJU�B�� �AY�p5��D.�O�U�`Վ�'a�b=��T� ]��\��BDIRa�i�� ��"��0DYN쒨���T�6 �R��,P&@���OPWOR�� ��,�@SYSB9U �SOP��c�$����U��� P ����PA����C2�+OP^`U�!��!xXB�AI�IMAGS�1�0U�7BIM��o��IN��@�n�RGO�VRD��	��K�P M�m�0� ߀�s��H2�L�B=з �PMGC_E�`cъANM��A�B1�BP��sSL�t�� ��0�OVSL�&S�D#EX�q}p/2G2� ��_��G�`��G�` Qfa�B�C�0p�%�c��_ZER�����s�� @hвb5O`RI��s0
��P�	��H��PL�Ĵ  _$FREE��E��Qq�!�Ls����yTD0;@ATUS㰎�AC_T��r�UB �_H��s�A4�`t�� D�AI�2RL��a2S�an S���XEY����1�� �0XUP��p��qPX�PF�D3����G�Ÿ��$SUBGb5��G��JMPWAIT8�V_%LOW�BQ��@CVF�QZPG2bb!Rz���U3CC� �R��MR�'IGNR�_PL�DBTB2;@P�qH1BW�P�$2��UP�%IG0�P=IG3TNLN�&2�R�����N�P)P�EED�8HADCOW;@�����E7pS4F1!4pSPDs�� L�0AV�5ps0�3UN�0"+0!R��LY�`� QNw��P��v1�G�C$��M�P�@L+.�NPA�T�2xDN��PIP%w0���ARSIZ�T��c�|q�Om`�h�AT�T���"\�B$�MEaM�B�A>C�3UX������`�ļ� $���SWIT�CHZ"�AW��ASr�8сCLLBv1��� $BArZ�D�s�BAM� h���I��@J50�����B6�F�A_KN�OW�3R��U!�A�D�H۠~0D��5YPAYLOA鱱�SS�_s�\W��\WZYSL�A�mpLCL_�� !���R�A����T���VF�YC�K��Z貓T��I�XR�M��W_ҬTB���JL)a_J�Q����AND^�9�8d�R�Q�w��PL�@AL_ ��@~0���A��k�C"�DXSE!��sJ3M`af� T���PDCK��r�C}OŰ_ALPHqc��cBE��W�qo�l��Т�!�� � ��40R_D_1YZ2�TDŰAR�4x!uxEv0s��TIA4_yu5_y6"�MOM��@ks�sxs�s�s��Bv �ADks�vxs�v�sPUB��R�t�uxs�uƅrk0�Ap��?� L$PI�1�s��^W.��xY.�I
:�IH�IV�<p}Q7��!�� !��b��8���73HIG�C73 w%p4Іp4w%� z�І��߈�!!w%SAMP���B�ЇC�w%�@>c 5�q��� 7 �Ҁ� ��p0"p�� 0p������hp���	���INќ�&�ؘ���ϔw"ښ���:�G�AMMƕS[%��$GET��o��D4�d��
ϡIB��2]I0�$HI�_��HsЩү�E�м�A��٠ʦLW�����٩@�ʦ�b��0caC�%GCHK��� 	��nI_%�����\bxΑ������s���v���c ��$�h 1����I� RCH_�D��'� �$)�LE@�������hذ�0_MSWFL�$M�`7SCR
(75_����3��dƧ���kp���x�p0�ĴDSVv1�P��v�Kǿ�	���S_SA�A�����NO�`C���d�� ��d_v_\�J�:ۂ�+R��w�0sD<�4��� 40��zʴ�ʈ��چ�1�����ՕәS/�@M��� � ��YL,�a������-� ��-���b��9�a�z�K����W�{� ���py�Ȳ�M� ���P��`a�$ 7���"�M���� �8 $���$W���ANG]�Q���d���d���d��d� נN�P���C��ϐX�0O��cΑZq��� ��[ �<�OM��"���1�C�U�g�bpCO�N��5L�a_�B� |�a�����y7xs 7�s��dzdO~z�AF�� B��ǲ@��PP-A�PM�ON_QUG� �� 8�0QCOUܴ�ǀQTH� HO�&�� HYSD@ES��B� UE� ��@O.5$�  �@P�৥N��RUNZY��09O��� � POP+�%���2ROGRQA���0:�2�Ov�+IT�xIN;FO��� �A_ğ8���`��� =(ʰSLEQ�����b�S_ED�d � � ���r�KԙQI#��EȠNU�'(AUT��%COPY�Q��8,����M��NB F+U�PRkUT� I"NF2U�B$G0�$��_RGADJ!�B3X_��2$�0�&~��&W�(P�(��&�73� �NH`_CY�C�	�!NSD9���LGOb����NYQ_FREQ��rW����^1RD)L��P:BV0�!�s���CcRE���c�IFH��jNAK�%�4_}G�STATU <å�MAILI�S�&@V��ǀLASTx�1�a04ELEM:1w� �EaNAB��0EASI&A��v� n�?�B���GF�����I���U2���� L�|BAB�C	PRS�LV	A�Fa�I���q1U����JP'c�F?RMS_TRvCΑ ��Ci����A�D��22��& 	SB 2�  �V�� 9V(b8WR��RNTdW&�
�DO�P�W}���04PR �;0��G�RID}�BAR�S��TY'C�ἐO\�p!� _�4�!� �R�TOo�74�� � |� PO�RXc�	bSRV��0)(d fDI��T�!pAaTd��^g��^g4�\i[�^g6\i7\i8�@a.1Fj�:1�$VALU�C��9D���F65�� !!"E��l�S�1��F_@AN���b�1R |c17ATOTALH�,�qCsPWK3I�QYtREGENWzlr��X�H@c5v� T1R�C�Wq_S���wlp\CV�!���u���1GRE�3�P�6B+�.  sV_H�PDA8���p�S_Y�i��o6SV�AR��2�� �"IG_SE��3�p b�5_/�tC=_�V$CMP���KDE�M���Ie��Z��^��� F�H�ANC�� p�&Q$E�2���IN�T?`iq��F%�M�ASK=��@OVR�3P� �P��1Α�Wp!��T� 4� �_XF�{�V�PSL9GV�:1� @K�� p5a���ApJpSh��4��U>�!���sTEa��`���`��U�Jd���3IL�_M~4���p� T�Q� ����@-�\�V�4�CB�P{�4AL�M�c�V1b�V1p�2��2p�3�3p�4�4p����p:����p���j�|�IN�VIAB��<�)���0�2,�U28�3,�38�4,��48� hR����� ��T $MC_YF�  ���L��(��ׅ7pM8�I׃����S ( ��n�K�EEP_HNADED��!ﴙ@��C��0��Q��?��O ��| ���p�܇�REM'��Iqb�L�c�h�U�4e�HPWD  ��SBM��PCOLLAB��p��5q�2��IT50`�w"N=O��FCAL�n�� ,��FL�>�A$SYN����M� Cq��XpUP�_DLY!�DGELA?�Jq�2Y� �AD���QSK;IP�� �`-�O;�NT�]�i�P_-V��^U�ip�� �q���q��u`�ڂ`�� �`�ڜ`�ک`�ڶ`��=9wA�J2R0� -�L�EX�@TX3N� �7AN� �N�}��4�RDC��� �:��Rz�TOR� ;���R�1�����;TR�GEA�rh@��RFcLG�^�5�ER����SPC�1UM�_N��2TH2N�1�A� 1ߏ ��A��Q62 � DKш��@O2_PC3]�S��|�1_0L10_C}2q 2��� �� $b� ���	V=� ����0�� �� S�b����mrj��CP��2��=��ID� �Gy�XUVL1a�1�n��� 10c�_D�S��=���1�Fv�11!� l�`����#C��ATE� �$�Q��bf���;T�3�HOME�� i2n��t����� �h3n���'9K 2f4n�n�����
]5n���/!/(3/E/]6n�h/z/��/�/�/�/�7n���/�/	??-??? 0��!8n�b?t?�?��?�?�?]S���!�  �Ag�p���Qc�Ed� T0C�tD:vtCIOꑔI�I@f�O��_OP��E�C4r��}�� WE�� ^@�l�q�P5�5s ����B$DSB��GNA��3s:�C��`���RS232zE� Ɍ���5���ICwEUS=sSPE(�>�aPARIT �2q�OPB���bFLO�WO�TR9@?rt�U�X�CUuP���aUX�T��a�ERFAiCZTT�U.pcwSCHa� t�b��_`Py���$ �&�pOM8���A�������UPDư��q3PTU@��EX��#hc�EFA8������RSP�P�a��|�`�7$USA�X��9��EX�PI��$(`�pY�eR_$�q�`mQ�fWR�OI�D���f��FFRI�END��L�$U�FRAMc�pTO;OLvMYH��r�LENGTH_V�TE�dI�;s��$Z pJxUFIN�V_^ ��_ARGuI%���ITI��bBwX�Sw�vG2�gG1�aꀎc�r�w�_r�O_XP��L�+q4���N�Sc��Cp�Pr�q��G���Rǁ󐒧�XQ؂��h�U���U��������PUd�X nm`E_MG`CT�c�H��h���U�dScG��W�`ć��لD]и@KȅJӂй�������$-� 2!���an �i1�h�`U2�k2=�3�k3�j -����iK���F�`l�P�`x�|�NtV�uV�ТPq,��r�P��� �V������R��pr�.���E9�<�Os�)E$A��T�P!Rh�U�k�ǓS��P���]Sb;Q� ! �ႃ"��K��"����S`�p�p��
��$$C��S��[��c ��9�9�� ؠVERSIܧ`���i��I#PP��AoAVM_�a2 �� ?0  �5�V�rb�S��� ��A	������9� �����ζ����ϧ�`�R�d�l�0�BS^ �r1�� <@ϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����|»CC`XLM�@v����  d��IN����qEX$?��2_`=�r ���0�IOCip,q ��PZXQ���{�IO'PV �1=�P $-��`ұ�!̺ �?�� � ��//%/7/I/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�o�o�o�o �o�o�o#5GY k}������ ���1�C�U�g�y� ��������ӏ���	� �-�?�Q�c�u����� ����ϟ����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i��{ύϟϱ���� LA�RMRECOV �I��LM_DG �����_IF ���p߂ߔߦ߀��^���������, 
 �G���@�m�����$_� ������ �2�D�V��h��NGTOL � I 	 A�   ����� PPINFO %� $������  1�I
�8 r\������� &W�p�Rd v��������//*/x�PPLI�CATION ?}����LR Ha�ndlingTo�ol y" 
V�9.10P/25���5'
8834�0z#�*F0�!�/1�31y#�,�/�"7�DF1� 5,y#No�ne5+FRA�5/ 6�-B&_�ACTIVE�� � [#��  X3U_TOMODb0)����U5CHGAPO�NL�? �3OUPLED 1M�� �0�?�?�?O;�CUREQ 1	�M�  TIL�L	XOiE_ ~D�wB�m%�MDH6E�2cJH�TTHKYwO��D\COUO_�O7O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q� c�u�����󏽏Ϗ� ����)�;�M�_�q� �����˟ݟ��� �%�7�I�[�m���� 믵�ǯٯ�����!� 3�E�W�i�{���翱� ÿտ�����/�A� S�e�wω��ϭϿ��� ������+�=�O�a� s߅��ߩ߻������߀��'�9�K�CET�O��d?X2DO_CLEAN�?V4���NM  �� O*�<�N�`�r�NDSPDRYR��&U5HI�0�@��� ��&8J\n�����R8MAX@I ��|�~A�7�X����!�2�!X2PLUG�G�0���3t5PRC*��B������.O3����SEGF�0Kz�������//&/^�LAP����Cz/�/�/ �/�/�/�/�/
??.?�@?R?�3TOTAL���3USENU
��; ��?~B@�RGDISPMM�C��AC��@I@���4O������3_STRING� 1
�;
�kM�0ST:
)A�_ITEM13F  nT=OOaOsO�O�O �O�O�O�O�O__'_�9_K_]_o_�_�_�_�I/O SIG�NAL-ETr�yout Mod�e4EInp�PS�imulated�8AOut�\�OVERR�� =� 1007BIn� cycl�U8A�Prog Abo�rc8A�TSta�tus6C	Hea�rtbeat2GMH Faulug~cAler�i�_�o �o�o�o�o $6H ��/K��AO K������� �)�;�M�_�q�����৏��ˏݏ_WOR �/K���=�O�a� s���������͟ߟ� ��'�9�K�]�o�����PO-Kia��-� ��ܯ� ��$�6�H� Z�l�~�������ƿؿ����� �2ϴ�DEV��]�ЯJτϖϨ� ����������&�8� J�\�n߀ߒߤ߶���>��PALTu}� -���)�;�M�_�q�� �������������%�7�I�[�m���GRI� /K�������� ��'9K]o �����������0Ru}I��# q������� //%/7/I/[/m//�/�/�/7PREG �� a�/?'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OGOYO�]��$ARG_�D ?	����A��  �	$�V	[��H]�G��W�I�@S�BN_CONFIQG�P�K�Q�RQ��ACII_SAVE  �TQS�@�TCELLSET�UP �J%  OME_IO�]��\%MOV_H8VPi_o_REPL�_��JUTOBACK�AQ�IQF�RA:\�+ X�_�&P'`T`�'�h� k
P �18/02�/09 11:0/6:04�&�H�-`{o�o�o�o�\���o�%7I[�&� �o������n ��+�=�O�a�s�� ������͏ߏ�|���'�9�K�]�o���X��  �Q_�S_\A�TBCKCTL.TM����ҟ����.�[INI�AeV~�SMESSAG!P�/�Q�@SQD�ODGE_D[P$VUb��O_�q��SPAUS�͠ !��K ,,		��@�Eѯ ߧů������Y� C�}�g�y�����׿���ӿ�������TSK  ��o��P�UPDTh�-�d�~�~�XWZD_E�NB-��J��STAp,��A~ŎAXIS�@?UNT 2�EQ�P� 	D���p��� &~��X���?�HF�*�� ��  X$U/k�>���-�  ����X;`UX��Tߍ�Pߊ�����ME�TK24�-S P���A�AK]�*A�{/6��1Ad�
A;�L��75n�8��S8cff4��DD7��6���@��SCRDC�FG 1�EN�Q �)UR�� ���������o�*Q%Ys�0�B�T�f�x� �������������,�����G�QGR`��r���k��NA�P��K	�Th_E�D+�1V�� 
� �%-��ED�T-Y�Z�M�D
TzP-�S��*�B��otV��  ��u2~�[\��� '�/Yk/�w3J/��/��s/�/ %/7/�/[/w4?�/ c?�/�??�?�/?�?'?w5�?R?/Ov?��OvO�?�?eO�?w6 �OO�OBO��OB_�O�O1_�Ow7z_�O�_ _��_oU_g_�_�_Bw8Fo��o���oo�o!o3o�oWow9�o_�o��;�`�o�o�#wCR} �_*�<��]�p����_��k � NO_D�E�yk GE_U�NUSEu�IG�ALLOW 1��	   (�*SYSTEM*���	$SERV�_GR��*���RE�G3�$U���*�N�UMX�}�k�PM}U�LAY�����PMPA�L,���CYC10ķ�ʞ�����UL�Swѭ�G�̒��5��L�?�BOXOR=I\�CUR_,�k��PMCNV���,�10����T4�DLI��%�G�	*�PROGRA2�?PG_MI���F��AL¥�����B�*�$FLU?I_RESUЗX�b����������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯�������H��k LAL_OUT� �T�WD_ABORѐ��j�O�ITR_RTN�  st��O�N�ONSTO� z�� b�CE_RIA3_I��z�������FCFG ��
��s}��_P}A9�GP 1����Q>�P�$b�!�C/�����z�-C�C ��(����+C8��@��H�� �CX��`��h��p���x}�����
�������	�su?���HE��O�NFI��Y�3G_mPr�1�� �� ă�}��������3KPAUSfI�1`�� �� �C`1oU� ������/5/@/Y/k/Q/�/Mo�NFO 1`��� � 	�-��//�� �"�D�A�/?������µ��B�QK��� D��b����B���B�3�0S��B��� 0²���B���j��r7�5B��a�80��O�����swV2LLECT_���&A���~7�EN z���2W1N[DE�3�7e����1234567890�7~rD����?�6ss
 ���q)9O^OD�8OJO�OE� |O�O�O�O�O�O/_�O __w_B_T_f_�_�_ �_�_o�_�_�_Ooo ,o>o�oboto�o�o�o��6B�2�; |�=�2IO  �9 �1yxy�as��/w�TR�2!}�� bJy
�o�~> ">}x�z���9_MORr#
� �'	X��!X� p�^���������1� �*q$?�,C?,,	��/�K�TqJr��%P[2&�?"�+�a�s�����
R���t7���u�y���5���s� ���9PDB�/�(7��dcpmidbg�]�v o�:��nD�pI���m�_  ��nG�毱��ï��.�����mg�x�C��Ůfg����-ſ�`ud1:���z'�?DEF 'y(Is�)��c�buf.txt�g��%��_MC8�)7�!sd�ō�7�*��������>|�Cz  B3A� �ClCy�C�d;�p������-D���D���D�J0?�M�D�I�D���~�-F����F��F�U��CH�S�F���*����,|P��t7A�pH �p�H �H ��t
����� E�@ Da�  D�  E	?� D�@ ��;��| Fp F�"� G=�fF��G'i�-�G>�Gg� �GK  H�<=�H�&HyM�c��  >�33O  `C/��n)���5YT娂��A��|�=L��<#�� �Vq����ξ��R�SMOFST �%8ʝ/P_T1���DE -3�c���q��Tq;�������?���<s�;��EST2�)+8�PR�2.a?��V��C4���|���p���������C��B͖��C�����H��p:d� ���T�_2�PROG ����%x�V$INUSER  �5�($KEY_TB�L  �"�	
��� !"�#$%&'()*�+,-./�7:;�<=>?@ABC�2�GHIJKLM�NOPQRSTU�VWXYZ[\]�^_`abcde�fghijklm�nopqrstu�vwxyz{|}�~���������������������������������������������������������������������߾����0���͓��������������������������������������������������?������q* �LCKt��&t S�TAT���_AU_TO_DO�6����IND�4�V1R����T27/�S�TO@/� TRL^, LETE�7~*�_SCREEN �?�kcs�c�2Uo MMEN�U 1/.� <ED?[�/?J? ճ'?M?�?]?o?�?�? �?�?�?�?O:OO#O pOGOYO�O}O�O�O�O �O�O$_�O_Z_1_C_ i_�_y_�_�_�_�_o �_�_oVo-o?o�oco uo�o�o�o�o
�o�o @)vM_�� �����*��� 9�r�I�[������ޏ ��Ǐ�&����\�3� E���i�{���ڟ��ß��Ϲ�#_MANU�ALs/�!DBCO� RIG�'�/�_oERRL2 0���a�N�����ǯ >P�NUMLI;�Z!�����
P�PXW�ORK 11�����'�9�K�]�o��D�BTB_�! 2���ç����D�B_AWAYX�^a�GCP ��=E�ö_AL;��òT��Yr �%��I�_r� �13#� , 
��T��B�ω�_M� I��Ѽ@����OoNTIM�'��������
�$�MOTNEN��z$��RECORD 1�9�� ��ψ�G�O�O�=߈�Ҳ{� �ߟ߱�Hع���O�� s�(�:�L����߂��� ��������� ���$� ��H���l�~������ ��5���Y� 2D ��h�������� �U
y�Rd v����?� //*/�N/9/G/�/ ��/�/�/;/�/�/q/ &?�/J?\?n??}?�? ?�?7?�?�?O�?�? FO�?jO�?�O�O�O�O _O�OWO_{O0_B_T_�f_�OòTOLER7ENCдB��ް�L��P�CSS_�CNSTCY 2�:����i_�� �_�_�_oo'o9oKo aooo�o�o�o�o�o�o��o�o#�TDEV�ICE 2;�[ ��vu��� �����*��ϭS�HNDGD <̼[�Cz|{�TLS 2=]}<������Џ����>��RPARAM >0�� |��}�SLAV�E ?]�I�_C�FG @J�*�d�MC:\�PL�%04d.CSV�)���cџ�RA &��CH�o�o�*�(�F��w�*�6�c��s�a�`��JP�Г�|����r�_C�RC_OUT �A]}��.�_NOC�OD~�B0���S�GN C&��&�j��21-�APR-21 0�0:38�*��09-FEB-18 11:06���v LIX��v�r�*�s�Iu5��M��Þ���������VE�RSION �-�V4.2.�10��EFLOG�IC 1D�[ 	��+�ɘ�!���PROG_ENqB�e�A�ULS��� d��_ACC�LIM���������WRSTJ�NT���*��MO�J�����INIT� E�Z&�*� ��OPTy� ?	�����
 	Rg575*�+�740ٕ61�71�5�[�1�U�21ԋ����TO  ݉����]V��DEX��d���p���PATH 9ۦ��A\��9��K�[HCP_CL?NTID ?Ѷ�� ��"S��Q�IAG_GRP {2J�� Q� 	 @K��@G�?����?l��>�������Q ������P)��?�b��?PT�i�^?տVm?Sݘ���f403 67�89012345�{������ ��s���@nȴ@i��#@d�/@_��w@Z~�@U�/@O�@I?��@D(������@���p����P�A�P�P�B4B��jp��ط�
���1��-@)h�s@$��@ bN@��@�����@�D@+�����������	 ��R��@N�@I�@D��@>�y@9@4� .v��@(��@"�\�Pbt��L��@Gl�@BJ@<z�@6��_0�`@*� $N�@���� $=q�@���F@�|�@33@��R@-?����?��`?��+hz�����Y"J�-@&��@N����!?�?� ��//*/</�- �/?�/&?8?�/?Z? �?^?�?�?@?R?�?�? O�?4OFO�?VO��ိ�9�Q�i @���V�AY����?��z��A��5AF��A4��@��L�4R��A��@��p� R�Q�R-�PP��@�� ��A�h��=H�9=����=�^5=��>P��>����=�,d_�,�P� ���C��<w(�U\� 4��l��_����A@��?��pO�_xM�_o0o �ȡT<ofo ovo�o~ox�o�o|I>��y�b��R=���=��zq���G�G��� � ��!�!�NUt@�T��V�쟷uB�� B��B��B�%�����~'����u���q�q6|��\�&���g���)PUB3pB�B A��@�"���m���<���  3���T�40�T�����g9y�f�wڔ�����D��\��3aB��Fp�l���r�ݏȏD��x�"�������3�����B���?�Ǐ p�돔������ܟ��9Q�0T<��I�;�������ν�XѶ�E�=����CT_CONF�IG K�m��eg7Ų�ST�BF_TTS��
@YɈ�Ȱ���������MAU��N�N�MS�W_CF\�L�� � ��OCVIE�W��M��ᄀ ��A�S�e�w������� /�Ŀֿ����ϭ� B�T�f�xϊϜ�+��� ��������,߻�P� b�t߆ߘߪ�9����� ����(��L�^�p� �����G����� � �$�6���Z�l�~���X����D�RC�N(E��!P�����!E�4iX���SBL�_FAULT �O����GPMS�K���P�TDIAOG P`��qo���o�UD1�: 6789012345t�n���P*�Sew�� �����//+/ =/O/a/s/2���R�
B�/J�TREC	P�
?)�+ A>?P?b?t?�?�?�? �?�?�?�?OO(O:O�LO^O�/�/�/�O�U�MP_OPTIO1N����ATR袒�:�	�EPME���O�Y_TEMP  �È�3B�r5P��TUNI͠���5QܦYN_BR�K Q��EDITOR�A�A_�R�_� ENT 1R���  ,&/MAIN��-�OdM?&PICK�_o� &DROP��_3o�PPROG_#o`o&}�os��to�o�o�o�o�o �o/SeL� p�������  �=�$�a�H�p���~� ����ߏ�؏����P�MGDI_STA�HU$�5Q}UNC;�1S� �dO��v�
�N
�Nd�Oݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W��En������� ��ʑ��ؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� ��g�q߃ߕߧ����� ������%�7�I�[� m����������� ���!�3�E�_�i�{� �������������� /ASew�� �����+ =W�Es����� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?Oak? }?�?E?��?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_G?Y?c_u_�_�_�? �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7Q_[ m��_���� ��!�3�E�W�i�{� ������ÏՏ���� �/�IS�e�w���� ����џ�����+� =�O�a�s��������� ͯ߯���'�A�3� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��9�K�U�g�yߋ� ������������	�� -�?�Q�c�u���� ������������C� M�_�q����ߧ����� ����%7I[ m������ �!;�EWi{ ��������/ ///A/S/e/w/�/�/ �/�/�/�/�/??3 !?O?a?s?��?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_+?=?G_Y_k_ !_�?�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	#_ 5_?Qcu�_�� ������)�;� M�_�q���������ˏ ݏ���-7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� %�/�A�S�e��q��� ����ѿ�����+� =�O�a�sυϗϩϻ� ���������9�K� ]�w����ߥ߷����� �����#�5�G�Y�k� }������������ �'�1�C�U�g��ߋ� ������������	 -?Qcu��� ����m��); M_y������ ��//%/7/I/[/ m//�/�/�/�/�/�/ �/!?3?E?W?q{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O?�O+_ =_O_i?__�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o__#5G�os_ }������� ��1�C�U�g�y��� ������ӏ��o� -�?�Q�ku������� ��ϟ����)�;� M�_�q���������˯ ݯ�	��%�7�I�c� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ��������� �/�A�[�M�w߉ߛ� �߿���������+� =�O�a�s����� ���������'�9�S� e�o������������� ����#5GYk }�������� 1C]�gy� ������	// -/?/Q/c/u/�/�/�/ �/�/I�??)?;? U_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�/ �O_!_3_M?W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�O�o+ E_;as���� �����'�9�K� ]�o���������ɏ�o� �$ENETM�ODE 1TFu��  
�`�`�e�"���RROR_PRO/G %��%�fe��r�@�TABLE  ��P��ß՟��@�SEV_NU�M �  ��	��@�_AU�TO_ENB  q,��=�_NO�� U��!���  *�]��]��]��]��+\�v���<��6�FLTR"�4��HIS��a�/�_�ALM 1V��� ��d]��`+ ��6�H�Z�l�~������_��<�  ���[�"�պ�TCP_�VER !��!�]���$EXTLO�G_REQ֦�-�'�SIZ0�"�SkTKM�K��$¿TOL  �aD�zޢ�A "�_BWD��������'�v��DI�� WFu��� ��a��S�TEP�������O�P_DOo���FD�R_GRP 1X����d 	пm�"��^�n&����c?��$,�MT� ��$ �����^ӳ����^�B��%BZ���B�S�B�?ȱB=�����(UB $B��V�Ae~�A��A����� ��:�%�^�I��m�����  AJAs�Y>(������`
 E�� x	����a?�{�������?�*�c���A�@����@�33@%�������@����L�����^�F@ ������������L��FZ!D�`��D�� BT��o@�����?���O��6���u���5�Zf5��ES������J��ƿ� .H�� ��X[x��n�4x�FEATUROE YFu��&��LR Ha�ndlingTo�ol ��bE�nglish D�ictionar}y�4D St� �ard��Analog I/O#�,gle Shi�ft?uto S�oftware �Updatedm�atic Bac�kup�	�gro�und Edit�� �Camera�:F>Commo�n calib �UI��n��M�onitor�t�r� Reliab<S�DHCP��
�Data Acq�uis�%)iag�nos�7?+oc�ument Vi�ewe"''ual� Check S�afety��hanced��
�%�s� Fr��xt�. DIO �f�iu$�'end� E�rr Lt"	=�'s�9r5�  ���
F�CTN Menu� v##[7TP I�nJ0facq5�G�igE�>�5�p �Mask Excھ g�'HT�0Pr?oxy Sv�$�6igh-Spe� �Ski��6m � m�munic�onsHurh0J0:/;��2connect� 2:Hncr�0sGtru8Ja@e�!� Jt%�KARE�L Cmd. L��0ua�8�CRunw-Ti� Env�H^K0el +�s��S/W�Lice�nse�#�,0Bo�ok(Syste�m)�
MACRO�s,�2/Offs	eZUH� w8/"P#MR �s.M}M@�!l�,MechStop�1tQ@Y"Ui2V�Vx� 7��L^odTwitc�h�_aSh!.BV�[O�ptmoaS�0fi�^aVg0GUult�i-T�0��	PC�M funkG�iaN�Ptiz~h�goV$/RegiPr@�f�ri� F�k�f8N?um Sel�U�i>�  Adju@�nx qV1}tatu�a�I�*�RDM R�obotsco3ve�ueav`� �Freq Anl�yGRem�P�!n��u�rServo�� �P�SNPX �b�B[SN�0Cl�i�!�WLibr�(��  �T:��voz�@th0ssag~e��� l5Q&�/�I�=��MILIB�����P Firmtu��Ph3Acc���TPTX4/��eln5PǏ���1U���orquTimu�la!�E�u�PPAa�A���!!c&�0gev.��mri� ��USR EV�NTğ֐nexc'ept� �pn�#ѕ,�(@VC�rBB�XVU 6��G�:�A��S�SC�y�SG�E����UI&Web Pl`vǮ�q0O���0�$�!?6ZDT� ApplD�
i�P0a!�:� Gr{id�qplay=�(���W�R-�.���h!N��B^P}200yiV4+scii�1�rLoad� �U�pl���f@I�Pat�V�ycS�B�`��� \6RL��� ۩~�5MI Dev�@� (�qR�f�?�gs�swo!�_64MB DRAMM����FRO�Ͼell:�sh��#בc.k �rp��5�t�ySs
r7̬r'`.�?+�p�!"=-o� 2z�a5port�.h�p�r q�-T1 ��{]P��No md�pc$筴OL���Sup��Fa�hOP�C-UA�l�T ȁ2eϓ�S0�0croa|�s:����~��Яuest�uS��eN2texV��up�1��#��PP�00�oV�irt�!�sR�st�dpnÛ�� SWIMEST f F0��������� �������� M DVpz���� ��
I@R lv������ ///E/</N/h/r/ �/�/�/�/�/�/?? ?A?8?J?d?n?�?�? �?�?�?�?O�?O=O 4OFO`OjO�O�O�O�O �O�O_�O_9_0_B_ \_f_�_�_�_�_�_�_ �_�_o5o,o>oXobo �o�o�o�o�o�o�o�o 1(:T^�� ������ �-� $�6�P�Z���~����� ��Ə����)� �2� L�V���z������� ����%��.�H�R� �v����������� ��!��*�D�N�{�r� ���������޿�� �&�@�J�w�nπϭ� �϶���������"� <�F�s�j�|ߩߠ߲� ���������8�B� o�f�x�������� �����4�>�k�b� t������������� 0:g^p� �����	  ,6cZl��� ���/�/(/2/ _/V/h/�/�/�/�/�/ �/?�/
?$?.?[?R? d?�?�?�?�?�?�?�? �?O O*OWONO`O�O �O�O�O�O�O�O�O_ _&_S_J_\_�_�_�_ �_�_�_�_�_�_o"o OoFoXo�o|o�o�o�o �o�o�o�oKB T�x����� ����G�>�P�}� t������������� ��C�:�L�y�p��� �������ܟ��� ?�6�H�u�l�~����� ���د���;�2� D�q�h�z�������ݿ Կ� �
�7�.�@�m� d�vϣϚϬ������� ���3�*�<�i�`�r� �ߖߨ���������� /�&�8�e�\�n��� ������������+�"� 4�a�X�j��������� ��������'0] Tf������ ��#,YPb �������� //(/U/L/^/�/�/ �/�/�/�/�/�/?? $?Q?H?Z?�?~?�?�? �?�?�?�?OO OMO DOVO�OzO�O�O�O�O �O�O_
__I_@_R_ _v_�_�_�_�_�_�_ oooEo<oNo{oro �o�o�o�o�o�o A8Jwn�� �������=� 4�F�s�j�|�����̍�  H5�51���2�R7�82�50�J6{14�ATUP��545�6�VC{AM�CUIF��28H�NRE�5�2;�R63�SC�H�DOCV��C�SU�869�0^�EIOCl�4���R69;�ESET�$�:�J7:�R68��MASK�PR�XYT�7�OCOB�3$������37�[J6
�53��He��LCH�OPLGz$�0O�MHCR ��S��MATk�MC�S#�0��55�MgDSW�B�OPB�GMPRC���s�0�PCMS�5J����l��s�51/�51{��0/�PRS�69�7�FRDG�FRE�Q�MCN�93��SNBAx�f�SHLB�M
ǀ����2�HTC#�TMsIL􈳖TPA˖oTPTX<�EL۶ĸ���8�����J9�5_�TUTC�UE�V�UEC�UF]RG�VCC��OǦwVIPG�CSCkƧCSGk���I�W�EB#�HTT#�R�6v���CG6�IG��IPGS\�RCvG�DGB�H75/��R7�Ry�R66�O�2O�R6�R5�5��4��5��D0u6�F�CLI3��.�CMS˖0�#�S[TY��TO7�7��t�_�ORSǦ���M��NOM˖OL��$���OPIs�SWEND�L��Sy��ETSsּ�S�CP�k�FVR˖IPNG�Gene�È6� H�Z�l�~��������� ������ 2DV hz������ �
.@Rdv �������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p������	  OH551��2�
oR782�50�	�J614�	ATU]P5456�	�VCAM�	CUI�F28lNREv�
52[R63��SCH�	DOCV��CSU�
869z0+EIOC��4R69[ES�ET<ZJ7ZR{68�
MASK�	�PRXY|7�
OCOL,3<X m3�*J653��H�,LCH�*OP�LG<0�*MHCuR�*SJ;MAT��MCS;0[+55�+MDSW�;�+OP�+MPR�*��,]0PCM{5K�X +X0�+51K5u1[L0KPRSK+�69�*FRDkFwREQ�
MCN�
{93SNBA�^�+SHLB�JM[t��<2HTC;�TMIL��TP�A*TPTX\ZEL�JX0�8
�
wJ95�TUT�*wUEVK*UEC�*wUFRkVCC+l�Ok:VIPkZCS�C�ZCSG��I��	WEB;HTTf;R6��\CG�k{IG�kIPGS�j�RCkZDG�+H7�5KR7:+RYLRk66�,2�*R6�WR55k|4�[5�{�D06+F�|CL9I�<JCMS*�pn;STY[kTO�kq7���ORSk:tx M�LNOM*�OL�;�0�OPI^�jSEND�
L:kSY�ETS�j {[�CP�FVR*I{PNkZGene� �R�d�v��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶��������� �"�4�F�X�j�|�� ������������� 0�B�T�f�x������� ��������,> Pbt�����}� STD�?LANG��	 '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_�ZRBT�OPT�N�_�_�_�_�_DPN�oo*o<o No`oro�o�o�o�o�o��o�oted ��>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|����������0�B�  �K�i�{��������Í99ʅ�$F�EAT_ADD �?	�����~��  	ǈ ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��� �����������&� 8�J�\�n��������� ��������"4F Xj|����� ��0BTf x������� //,/>/P/b/t/�/ �/�/�/�/�/�/?? (?:?L?^?p?�?�?�? �?�?�?�? OO$O6O HOZOlO~O�O�O�O�O��O�O�DEMO �Y��   ǈ1]'_9_f_]_o_ �_�_�_�_�_�_�_�_ ,o#o5oboYoko�o�o �o�o�o�o�o�o( 1^Ug���� ����$��-�Z� Q�c�������Ə��Ϗ �� ��)�V�M�_� ��������˟�� ��%�R�I�[���� ������ǯ���� !�N�E�W���{����� ��ÿݿ����J� A�Sπ�wω϶ϭϿ� �������F�=�O� |�s߅߲ߩ߻����� ���B�9�K�x�o� ������������ �>�5�G�t�k�}��� ����������: 1Cpgy��� �� �	6-? lcu����� ��/2/)/;/h/_/ q/�/�/�/�/�/�/�/ ?.?%?7?d?[?m?�? �?�?�?�?�?�?�?*O !O3O`OWOiO�O�O�O �O�O�O�O�O&__/_ \_S_e_�_�_�_�_�_ �_�_�_"oo+oXoOo ao�o�o�o�o�o�o�o �o'TK]� �������� �#�P�G�Y���}��� ������׏���� L�C�U���y������� ܟӟ��	��H�?� Q�~�u�������دϯ ����D�;�M�z� q�������Կ˿ݿ
� ��@�7�I�v�m�� �ϣ����������� <�3�E�r�i�{ߕߟ� ����������8�/� A�n�e�w������ �������4�+�=�j� a�s������������� ��0'9f]o �������� ,#5bYk�� ������(// 1/^/U/g/�/�/�/�/ �/�/�/�/$??-?Z? Q?c?}?�?�?�?�?�? �?�? OO)OVOMO_O yO�O�O�O�O�O�O�O __%_R_I_[_u__ �_�_�_�_�_�_oo !oNoEoWoqo{o�o�o �o�o�o�oJ ASmw���� �����F�=�O� i�s�������֏͏ߏ ���B�9�K�e�o� ������ҟɟ۟��� �>�5�G�a�k����� ��ίůׯ����:� 1�C�]�g�������ʿ ��ӿ ���	�6�-�?� Y�cϐχϙ��Ͻ��� �����2�)�;�U�_� �߃ߕ��߹������� �.�%�7�Q�[��� ������������*� !�3�M�W���{����� ����������&/ IS�w���� ���"+EO |s������ �//'/A/K/x/o/ �/�/�/�/�/�/�/? ?#?=?G?t?k?}?�? �?�?�?�?�?OOO 9OCOpOgOyO�O�O�O �O�O�O_	__5_?_ l_c_u_�_�_�_�_�_ �_ooo1o;oho_o qo�o�o�o�o�o�o
 -7d[m� �������� )�3�`�W�i������� ̏ÏՏ����%�/� \�S�e�������ȟ�� џ�����!�+�X�O� a�������į��ͯ�� ���'�T�K�]��� ��������ɿ����� �#�P�G�Yφ�}Ϗ���ϳ��������  �+�=�O�a� s߅ߗߩ߻������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}����� ����������1 CUgy���� ���	-?Q cu������ �//)/;/M/_/q/ �/�/�/�/�/�/�/? ?%?7?I?[?m??�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao so�o�o�o�o�o�o�o '9K]o� �������� #�5�G�Y�k�}����� ��ŏ׏�����1� C�U�g�y��������� ӟ���	��-�?�Q� c�u���������ϯ� ���)�;�M�_�q� ��������˿ݿ�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w������� ������+�=�O�a� s��������������� '9K]o� ������� #5GYk}�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?u?�?�?�?�?�?�? �?OO)O;OMO_OqO �O�O�O�O�O�O�O_>Y  XQ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9K] o������� ��#�5�G�Y�k�}� ������ŏ׏���� �1�C�U�g�y����� ����ӟ���	��-� ?�Q�c�u��������� ϯ����)�;�M� _�q���������˿ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߱����������� /�A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?�?�?�?�?�?�?O O1OCOUOgOyO�O�O��O�O�O�O�O	_QPX3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ��� ������%�7�I�[� m�ߑߣߵ������� ���!�3�E�W�i�{� ������������� �/�A�S�e�w����� ����������+ =Oas���� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ �������� �/�A�S�e�w����� ����я�����+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ ����#�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	����$FEAT_D�EMOIN  V ԀK�� �3�_INDEX@�O���3�ILECOM�P Z������N�.�w�S�ETUP2 [������  �N ��t�_AP2�BCK 1\��  �)�����%��� ����H� ���t���'���� ]�����(���L��� p������5�����k�  ��$��1Z��~ ��C�g� �2�Vh�� �?��u
/�./ @/�d/��/�/)/�/ M/�/�/�/?�/<?�/ I?r??�?%?�?�?[? �??O&O�?JO�?nO �OO�O3O�OWO�O�O �O"_�OF_X_�O|__ �_�_A_�_e_�_o�_ 0o�_To�_ao�oo�o =o�o�oso�o,> �ob�o��'�K@�o������P��� 2��*.V1R�g��p*j���`�s�����uQ�PC|��pFR6:֏"���;�ʋT_�_� q� �\���B�,����v�*.FT���q	�������C�қSTM c�l�w��d�����piPen�dant Panel��қH�������该�3�L�ӚGIF V�����l�)�;�пӚJPGڿϋ�𿭿��T�ˊJS^χ��p��u�2�%
Ja�vaScript��޿CS��ߊ������ %Casc�ading St�yle Shee�ts7ߩp
ARGNAME.DTf�
�|��\z�8ߚ������g���DISP*�ߔߎ���>���0��?���	PANEL15��%��������ǯu�2����������o�z�3;����� ��L�^���z�4��%�������wr�TP�EINS.XML�~�:\�PbC�ustom To�olbar���PASSWORDC~�~FRS:\�� %Pass�word Con�figW��4�/ �ԝ[U�/qֱ䘯 ���/�b_/v���/%J(�/g/y/?'2T/=?H(+?�/�/ �?��?�/U5�?o?�?O'3\?EOH(3O�? O�O���O�?]E�OwO�O_'4dOM_H(;_ �O_�_�_�OeU�_ _�_&o�Jo�no� ��o3o�oWo�o�o�o "�oFX�o|� �A�e���0� �T��M������=� ҏ�s����,�>�͏ b�񏆟�'���K��� o�ٟ���:�ɟ^�p� ����#���ʯY��}� �����H�ׯl���e� ��1�ƿU������ � ��D�V��z�	Ϟ�-� ?���c��χ���.߽� R���v߈�߬�;��� ��q���*����`� �߄��}��I���m� ����8���\�n��� ��!���E�W���{� ��	F��j���� /�S���� B��x�+���a�,�$FI�LE_DGBCK� 1\������ <� �)
SUMM?ARY.DG/�]�MD::/z/��Diag Sum�mary{/([CONSLOGp/S/e!��/�/�!Console log�/~�\TPACCN�/�Y?%A?~?�%TP� Account�in ?�Y@6:I�PKDMP.ZI	P�?�
�?O�%�0�ExceptionO�*�_\O��bQJO�_1FR �DT Files��O�<f MEMCH�ECKt?�/i/_�1Memory �Data_�
l�)	FTP�/�f_�Oj_W1mm�e`TBD�_�L� >I)ETHERNET�_��A��_o�!Ethe�rnet 0fi�gura&O�}QDCSVRF�_m__ܘoQ%]` v�erify alyl�o�M.cXeDIFF�ovo�o� P%�hdif�f�g�A]`CHG01�o��a5,��b- `y2�@�&�1��gr3�8���� <�я�`�VTRNDIAG.LS֏�����.�!Q� Ope�>c Log �!n�ostic����)VDEV�DA}O�����a�VisQ�Dev�iceX�e�IMG@��?����4�7�ʔ�Imag֟c�U�P{�ESz��F�RS:\z��O@U�pdates L�ist���"�FLEXEVENo��%�>��a� UIF Ev�QU�?��  ,�sz)
�PSRBWLD.CMj���������0PS_ROBO�WEL�_�*�HADOW4��+�D��SShadow? Chang�O���a��RCMERR<�!�3���S���CFG Er�rorАtail>k� =��B��SGLIB�ϧϹ�tN�!Q� St?`x_�����):ЃZDU_��7���W�ZDT�adn����NOTIbo�߽��R�UNotif�ic?b��t��AGXbGIGE��/�A�<��]�GigEZ�d��N�A��-�� Q��^������:��� ��p���);��_ ����$�H�l ��7�[m� � ��V�z/ !/�E/�i/�v/�/ ./�/R/�/�/�/?�/ A?S?�/w??�?�?<? �?`?�?�?O+O�?OO �?sO�OO�O8O�O�O nO_�O'_9_�O]_�O �__�_�_F_�_j_�_ o�_5o�_Yoko�_�o o�o�oTo�oxo�o C�og�o��, �P�����?� Q��u����(���Ϗ ^�󏂏�)���M�܏ q������6�˟ݟl� ���%���2�[��� �����D�ٯh���� ��3�¯W�i������ ��@����v�Ϛ�/� A�пe����ϛ�*Ͽ� N����τ�ߨ�=��� J�s�ߗ�&߻���\� �߀��'��K���o� ����4���X����� ��#���G�Y���}�� ����B���f����� 1��U��b���>��t	�$�FILE_FRS�PRT  ���� ����$MDONLY� 1\8�  
 ��{��� �����///� S/�w/�//�/</�/ �/r/?�/+?�/8?a? �/�??�?�?J?�?n? OO�?9O�?]OoO�? �O"O�OFO�O�O|O_ �O5_G_�Ok_�O�_�_ 0_�_T_�_�_�_o�_�Co�_Poyo"VIS�BCKV@e*�.VD�o�o8`F�R:\�`ION\�DATA\�oZb�8`Vision� VD file �oo>Pfot^o� '��]���(� �L��p�����5� ʏ܏�� ���$���5� Z��~������C�؟ g�������2���V�h� #������?����u� 
���.�@�ϯd�󯈿��)���LUI_�CONFIG �]8�aɻ '$ ��[{8 π2�D�V�h�zψ��|x������������
� ��-�?�Q�c�u�߆� �߽������ߊ��)� ;�M�_�q����� ��������%�7�I� [�m������������ ����!3EWi  ������~ /ASe�� ����h�// +/=/O/�s/�/�/�/ �/�/d/�/??'?9? K?�/o?�?�?�?�?�? `?�?�?O#O5OGO�? kO}O�O�O�O�O\O�O �O__1_C_�Og_y_ �_�_�_�_X_�_�_	o o-o�_>ocouo�o�o �oBo�o�o�o) �oM_q���> �����%��I� [�m������:�Ǐُ ����!���E�W�i� {�����6�ß՟��� ����A�S�e�w���  �����ѯ������ +�=�O�a�s������ ��Ϳ߿�Ϛ�'�9� K�]�oρ�ϥϷ��� �����ϖ�#�5�G�Y� k�}�ߡ߳������� �ߎ��1�C�U�g�y��	���x����$�FLUI_DAT�A ^���>�����RESULT 2�_���� ��T�/wiza�rd/guide�d/steps/?Expert��"� 4�F�X�j�|���������������Con�tinue wi�th G��ance��1CUgy������� ��-����0� ������$���ps�o�� ������/#/ 5/���\/n/�/�/�/ �/�/�/�/�/?"?4?�F>$(:Jrip�X�?�?�?�? OO*O<ONO`OrO�O C/�O�O�O�O�O__ &_8_J_\_n_�_�_Q?�c?�_�?EJ�T�imeUS/DST�_"o4oFoXojo|o��o�o�o�o�o��Enabl
. @Rdv�������� �_��_�_f24or��� ������̏ޏ���� &��o�o\�n������� ��ȟڟ����"�4�����)�;�M�zon
`7�ʯܯ� ���$�6�H�Z�l�~����EST Ea�rn Stand�� ����ӿ���	��-��?�Q�c�uχ�� ��t�f�x�:���acces�?�+� =�O�a�s߅ߗߩ߻��������nect� to Network���%�7�I� [�m���������
�ȘA��Ϻ��ϊ��!��`Introduction�� t��������������� (�OL^p� ������ $5�_�P*���~�VEditor5 ����
//./@/�R/d/v/5 Tou�ch Panel� � (reco/mmen�P)�/�/ �/�/�/?#?5?G?Y?k?}?�̬P�^�?� B�?OO/OAOSOeO wO�O�O�O�O�O<�O __+_=_O_a_s_�_ �_�_�_�_�Y�0�?�:�?o�?EoWoio {o�o�o�o�o�o�o�o �OASew� �������� +��_�_op�2o���� ��͏ߏ���'�9� K�]�o�.������ɟ ۟����#�5�G�Y� k�}�<���`�¯��� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ��ώ��ϲ��֯ ;�M�_�q߃ߕߧ߹� ��������%��I� [�m��������� �����!���B��f� (�*������������� /ASew6� ������ +=Oas2��V� ����//'/9/ K/]/o/�/�/�/�/�/ ��/�/?#?5?G?Y? k?}?�?�?�?�?�� ��?O�COUOgOyO �O�O�O�O�O�O�O	_ _�/?_Q_c_u_�_�_ �_�_�_�_�_oo�?  O�?Dono0O�o�o�o �o�o�o%7I [m,_����� ���!�3�E�W�i� (o:oLo^o���o��� ��/�A�S�e�w��� ������~����� +�=�O�a�s������� ��ͯ�������ԏ9� K�]�o���������ɿ ۿ����П5�G�Y� k�}Ϗϡϳ������� ����ޯ��d�&� �ߝ߯���������	� �-�?�Q�c�"�t�� �����������)� ;�M�_�q�0ߒ�T߶� x�����%7I [m������ ��!3EWi {��������� /��//A/S/e/w/�/ �/�/�/�/�/�/?? �=?O?a?s?�?�?�? �?�?�?�?OO�6O �ZO/O�O�O�O�O �O�O�O_#_5_G_Y_ k_*?�_�_�_�_�_�_ �_oo1oCoUogo&O �oJO�o�o�_�o�o	 -?Qcu�� ��|_����)� ;�M�_�q��������� xo�o�o���o7�I� [�m��������ǟٟ �����3�E�W�i� {�������ïկ��� �ʏ��8�b�$��� ������ѿ����� +�=�O�a� ��ϗϩ� ����������'�9� K�]��.�@�R���v� �������#�5�G�Y� k�}����r����� ����1�C�U�g�y� ���������ߒߤ� ��-?Qcu�� �������) ;M_q���� ���//������ X//�/�/�/�/�/ �/�/?!?3?E?W? h?�?�?�?�?�?�?�? OO/OAOSOeO$/�O H/�Ol/�O�O�O__ +_=_O_a_s_�_�_�_ �_�O�_�_oo'o9o Ko]ooo�o�o�o�ovO �o�O�o�O#5GY k}������ ���_1�C�U�g�y� ��������ӏ���	� �o*��oN������ ����ϟ����)� ;�M�_���������� ˯ݯ���%�7�I� [��|�>�����v�ٿ ����!�3�E�W�i� {ύϟϱ�p������� ��/�A�S�e�w߉� �߭�l��������ƿ +�=�O�a�s���� �����������'�9� K�]�o����������� �����������,V �}������ �1CU�y �������	/ /-/?/Q/"4F �/j�/�/�/??)? ;?M?_?q?�?�?�?f �?�?�?OO%O7OIO [OmOO�O�O�Ot/�/ �/�O�/!_3_E_W_i_ {_�_�_�_�_�_�_�_ �?o/oAoSoeowo�o �o�o�o�o�o�o�O �O�OL_s��� ������'�9� K�
o\���������ɏ ۏ����#�5�G�Y� z�<��`şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u����� ��j�̿��𿲟�)� ;�M�_�qσϕϧϹ� ���������%�7�I� [�m�ߑߣߵ����� ���߼���B��� {������������ ��/�A�S��w��� ������������ +=O�p2�� j����'9 K]o���d�� ���/#/5/G/Y/ k/}/�/�/`���/ �/�?1?C?U?g?y? �?�?�?�?�?�?�?� O-O?OQOcOuO�O�O �O�O�O�O�O�/�/�/  _J_?q_�_�_�_�_ �_�_�_oo%o7oIo Omoo�o�o�o�o�o �o�o!3E__ (_:_�^_���� ��/�A�S�e�w��� ��Zo��я����� +�=�O�a�s������� hz��'�9� K�]�o���������ɯ ۯ���#�5�G�Y� k�}�������ſ׿� ����̟ޟ@��g�y� �ϝϯ���������	� �-�?���P�u߇ߙ� �߽���������)� ;�M��n�0ϒ�TϹ� ��������%�7�I� [�m������������ ����!3EWi {��^������� /ASew� ��������/ +/=/O/a/s/�/�/�/ �/�/�/�/�?�6? ��/o?�?�?�?�?�? �?�?�?O#O5OGO/ kO}O�O�O�O�O�O�O �O__1_C_?d_&? �_�_^O�_�_�_�_	o o-o?oQocouo�o�o XO�o�o�o�o) ;M_q��T_�_ x_���_�%�7�I� [�m��������Ǐُ 돪o�!�3�E�W�i� {�������ß՟矦 ���>� �e�w��� ������ѯ����� +�=���a�s������� ��Ϳ߿���'�9� ��
��.���R����� �������#�5�G�Y� k�}ߏ�N��������� ����1�C�U�g�y� ���\�nπ����	� �-�?�Q�c�u����� ����������) ;M_q���� ���������4�� [m����� ��/!/3/��D/i/ {/�/�/�/�/�/�/�/ ??/?A? b?$�? H�?�?�?�?�?OO +O=OOOaOsO�O�O�? �O�O�O�O__'_9_ K_]_o_�_�_R?�_v? �_�?�_o#o5oGoYo ko}o�o�o�o�o�o�o �O1CUgy �������_� �_*��_�c�u����� ����Ϗ����)� ;��o_�q��������� ˟ݟ���%�7�� X��|���R���ǯٯ ����!�3�E�W�i� {���L���ÿտ��� ��/�A�S�e�wω� H���l����Ϣ��� +�=�O�a�s߅ߗߩ� �����ߞ���'�9� K�]�o������� ����Ͼ��2���Y� k�}������������� ��1��Ugy �������	 -�����"��F� �����//)/ ;/M/_/q/�/B�/�/ �/�/�/??%?7?I? [?m??�?Pbt�? ��?O!O3OEOWOiO {O�O�O�O�O�O�/�O __/_A_S_e_w_�_ �_�_�_�_�_�?�?�? (o�?Ooaoso�o�o�o �o�o�o�o'�O 8]o����� ����#�5��_V� oz�<o����ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u���F� ��j�̯�����)� ;�M�_�q��������� ˿ݿ����%�7�I� [�m�ϑϣϵ����� ���ϼ�����W�i� {ߍߟ߱��������� ��/��S�e�w�� ������������ +���L��p���F�� ��������'9 K]o�@��� ���#5GY k}<���`����� �//1/C/U/g/y/ �/�/�/�/�/��/	? ?-???Q?c?u?�?�? �?�?�?����?&O �MO_OqO�O�O�O�O �O�O�O__%_�/I_ [_m__�_�_�_�_�_ �_�_o!o�?�?OO xo:O�o�o�o�o�o�o /ASew6_ �������� +�=�O�a�s���DoVo hoʏ�o���'�9� K�]�o���������ɟ �����#�5�G�Y� k�}�������ůׯ�� �����ޏC�U�g�y� ��������ӿ���	� �ڟ,�Q�c�uχϙ� �Ͻ���������)� �J��n�0��ߧ߹� ��������%�7�I� [�m��ߣ������ �����!�3�E�W�i� {�:ߜ�^��������� /ASew� ������� +=Oas��� �������/��� K/]/o/�/�/�/�/�/ �/�/�/?#?�G?Y? k?}?�?�?�?�?�?�? �?OO�@O/dOvO :?�O�O�O�O�O�O	_ _-_?_Q_c_u_4?�_ �_�_�_�_�_oo)o ;oMo_oqo0OzOTO�o �o�O�o%7I [m�����_ ���!�3�E�W�i� {�������Ï�o�o�o ����oA�S�e�w��� ������џ����� �=�O�a�s������� ��ͯ߯���ԏ� ��
�l�.�������ɿ ۿ����#�5�G�Y� k�*��ϡϳ������� ����1�C�U�g�y� 8�J�\��߀�����	� �-�?�Q�c�u��� ���|�������)� ;�M�_�q��������� ���ߜ߮���7I [m����� ���� EWi {������� //��>/ b/$�/ �/�/�/�/�/�/?? +?=?O?a?s?�/�?�? �?�?�?�?OO'O9O KO]OoO./�OR/�Ov/ �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�?�_ �_oo1oCoUogoyo �o�o�o�o�O�o�O �O�o?Qcu�� ��������_ ;�M�_�q��������� ˏݏ����o4��o X�j�.�������ǟٟ ����!�3�E�W�i� (�������ïկ��� ��/�A�S�e�$�n� H�����~������ +�=�O�a�sυϗϩ� ��z�������'�9� K�]�o߁ߓߥ߷�v� �������п5�G�Y� k�}���������� �����1�C�U�g�y� ��������������	 ��������`"�� �����) ;M_����� ���//%/7/I/ [/m/,>P�/t�/ �/�/?!?3?E?W?i? {?�?�?�?p�?�?�? OO/OAOSOeOwO�O �O�O�O~/�/�/_�/ +_=_O_a_s_�_�_�_ �_�_�_�_o�?o9o Ko]ooo�o�o�o�o�o �o�o�o�O2�OV _}������ ���1�C�U�g�x ��������ӏ���	� �-�?�Q�c�"��F ��jϟ����)� ;�M�_�q��������� x�ݯ���%�7�I� [�m��������t�ֿ ��������3�E�W�i� {ύϟϱ��������� �ʯ/�A�S�e�w߉� �߭߿��������ƿ (��L�^�"߅��� ����������'�9� K�]�߁��������� ������#5GY �b�<��r��� �1CUgy ���n����	/ /-/?/Q/c/u/�/�/ �/j���/?�)? ;?M?_?q?�?�?�?�? �?�?�?O�%O7OIO [OmOO�O�O�O�O�O �O�O�/�/�/�/T_? {_�_�_�_�_�_�_�_ oo/oAoSoOwo�o �o�o�o�o�o�o +=Oa _2_D_� h_�����'�9� K�]�o�������doɏ ۏ����#�5�G�Y� k�}�������r�� ����1�C�U�g�y� ��������ӯ����� �-�?�Q�c�u����� ����Ͽ���ğ&� �J��qσϕϧϹ� ��������%�7�I� [�l�ߑߣߵ����� �����!�3�E�W�� x�:Ϝ�^��������� ��/�A�S�e�w��� ����l������� +=Oas��� h�������'9 K]o����� �����#/5/G/Y/ k/}/�/�/�/�/�/�/ �/�?�@?R?/y? �?�?�?�?�?�?�?	O O-O?OQO/uO�O�O �O�O�O�O�O__)_ ;_M_?V?0?z_�_f? �_�_�_oo%o7oIo [omoo�o�obO�o�o �o�o!3EWi {��^_�_�_�� �_�/�A�S�e�w��� ������я����o� +�=�O�a�s������� ��͟ߟ���� H�
�o���������ɯ ۯ����#�5�G�� k�}�������ſ׿� ����1�C�U��&� 8���\���������	� �-�?�Q�c�u߇ߙ� X�����������)� ;�M�_�q����f� xϊ�����%�7�I� [�m������������ ������!3EWi {������� ����> �ew� ������// +/=/O/`s/�/�/�/ �/�/�/�/??'?9? K?
l?.�?R�?�? �?�?�?O#O5OGOYO kO}O�O�O`/�O�O�O �O__1_C_U_g_y_ �_�_\?�_�?�_�?�_ o-o?oQocouo�o�o �o�o�o�o�o�O) ;M_q���� ����_��_4�F� 
m��������Ǐُ ����!�3�E�i� {�������ß՟��� ��/�A� �J�$�n� ��Z���ѯ����� +�=�O�a�s�����V� ��Ϳ߿���'�9� K�]�oρϓ�R���v� ���Ϭ��#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ����������϶� ����<���c�u����� ����������) ;��_q���� ���%7I ��,��P���� ��/!/3/E/W/i/ {/�/L�/�/�/�/�/ ??/?A?S?e?w?�? �?Zl~�?�OO +O=OOOaOsO�O�O�O �O�O�O�/�O_'_9_ K_]_o_�_�_�_�_�_ �_�_�?o�?2o�?Yo ko}o�o�o�o�o�o�o �o1CTogy �������	� �-�?��_`�"o��Fo ����Ϗ����)� ;�M�_�q�����T�� ˟ݟ���%�7�I� [�m����P���t�֯ �����!�3�E�W�i� {�������ÿտ翦� ��/�A�S�e�wω� �ϭϿ����Ϣ��Ư (�:���a�s߅ߗߩ� ����������'�9� ��]�o������� �������#�5���>� �b���N߳������� ��1CUgy �J�����	 -?Qcu�F� ��j�����//)/ ;/M/_/q/�/�/�/�/ �/�/�??%?7?I? [?m??�?�?�?�?�? ����0O�WOiO {O�O�O�O�O�O�O�O __/_�/S_e_w_�_ �_�_�_�_�_�_oo +o=o�?O O�oDO�o �o�o�o�o'9 K]o�@_��� ����#�5�G�Y� k�}���No`oroԏ���$FMR2_G�RP 1`���� �C�4  B��p	 ��p�0��F;@ F�E��Q�F����C��L�FZ�!D�`�D��� BT��@��=�^�?�  ������6������5�Zf5�EySΑ^�A�  ����BH��\��@�/33@�� ���!�@�Q��@�g��]�Q����<�z��<�ڔ=7��<�
;;�*��<��^�8ۧ��9k'V8���8���7ג	8(��~���� �=�(�a�L����w�_CFG a��T0���ӿ�����N�O �
F�0+� 0���RM_�CHKTYP  ��p	�����R{OMF�_MINL���s��x��7�X��SSB��b��? �����u�����ϝ�TP_�DEF_OW  ��t	���IRC�OMK����$GE�NOVRD_DOrm��q*�THRm�� dG�d0�_EN�B� 0�RAV�C��c���� ��>�����v���^�����.� ��OUU��i�3�.��.�<u������,�z����sC� � D����l��$�@��B�/��1�m�\�ϑ�SMT��j���������$HOS�TC��1k���s��� MC�t�����v _ 27.0 1��  e��BTf x�
0�������	anonymous4FX@j|�r����� ����)
//./@/ R/�v/�/�/�/�i/ �/??*?<?N?� ���?�/�?��?�? OO�/�?JO\OnO�O �?�O�/�O�O�O�O_ S?�Ow?�?j_�O�?�_ �_�_�_�_+Ooo0o BoTow_�O�O�o�o�o �o�o'_9_K_]__o5 �_t�����_� ���(�K}o�op� ���������o1 3�$�gH�Z�l�~��� ���Ɵ؟����Q� �D�V�h�z���Ϗ� 󏥯���;��.�@� R�d������������ �%���*�<�N�`� ����ǯ��ۿ����� ��&�i�J�\�n߀� �ߵ�7�����������"�o���ENT 1�l���  P!\��s�  u�a� ���������
��� ���?�d�'���K��� o�����������*�� Nr5�Yk� ����8�1 n]�U�y�� ��/4/�X//|/ ?/�/c/�/�/�/�/�/�?�/B?:QUICC0O?+?=?�?a4A1�?{?�?�?a42�?��?�?>O!ROU�TER?OO-O�O!?PCJOG�OjO�!192.168.0.10h?~]3CAMPRT�O�O!�E1�@_�F�RTXO
__}_C�N�AME !P�!�ROBO�O�_S_CFG 1kP�� �A�uto-star�ted��FTP��a�Ϧ�Ao��eo wo�o�o�oF��o�o�o *o�oOas� ��r��_oo�' Io�<�N�`�r�5�� ����̏ޏ����&� 8�J�\�n�g�yϋϝ� 鏿�����"�4�F� 	�j�|�������՟W� �����0�B����� ���������ҿ��� ��ݯ>�P�b�tφ� ��+ϼ��������� Y�k�}�/ߑς�ſ�� �������߱��$�6� H�k�l��ߐ����� ����-�?�Q�2�e�V� ��z�������s����� ��
?���;dv �������%� 9[�<N`r�G ������&/ 8/J/\/n/�/��� ���//?"?4?F? X?/|?�?�?�?�?�/ i?�?OO0OBOTO�Z_ERR m�Z�\OlFPDUSIZW  �0^0��D�>�EWRD ?��U�!�  guest�6��O�O __$_6_�TS�CD_GROUP� 3n�\ �Q��9IFT|^$PA�|^OMP|^ n|^_SH|^ED�_w $C|^COMn@�TTP_AUTH� 1o{K <!�iPendan�BWMn�[�2�q!KAREL:*MoVohmKC}o�o�o�u`VISION SETfP�o�o�v!,rcP>h b������~dCTRL p{M�6��1
F�F�FF9E3��$�FRS:DEFA�ULT[�FA�NUC Web ?Server[�I� �"d�O�D�я������+�jDWR_C�ONFIG q.kU�Bc[�lA�IDL_CPU_kPCz��1B��  BH��MIN���sQ��GNR_I�OuA�B�0�H��NP�T_SIM_DO�ӖݛSTAL_oSCRNӖ �ޚ�TPMODNTOqL�ݛ��RTY��p����` `ENB��sS��OLNK 1r{KxP����ɯ�ۯ������MAS�TEҐy�5���SLAVE s{K�H D��SRAMCACHE/�A�"aO_CFGq������UO�`����CMT�_OPz�ՒJǳY�CLp���t�_AS�G 1t`��A
 �6�H�Z�l�~ϐ� �ϴ���������� �\�	�NUM�CI�
��IPn���RTRY_CNҿ���G_UP_��A����E� ������u)� � 06��م�RC�A_ACC 2v�k[  R��� �� �� 5� 7Þ��0i��,�. � p#��  ��2D���BUF00�1 2wk[= ��u��u0�Z���������#��2��C��Vu�0% Pou�0Bx2��u0�q��������u0�sWP���Ц�������2p  2�p�J��U.�c�u0�r`�|�u0Z�p���.��.��.��.���.��.�Ԗ�So2ݠ(�S�~��u�0!�SpS�u0X]�S�~���~��u0�p��S���T�q�  �qT ��/���@��d�  ��Tz���U�����������������QR��=��r�䃖�Y���]����Ö��s�2���d�� �����������������t�� ���tp ���t� x���� ���������%�&�,�``�4��<�AE�A M�AU�A]�Ae�A m�Au�A}������e ���� ��������������������W�������������U� (�����kX	�" � �x ���	l,p>Pbt003� �� ���1���" ����"����"��" ��"����"��"� �"�#�"%�3:2 5�C:2E�:2M�[:2 ]�k:2m�{:2}� �2����2��2�� ��2��2����2�� �����2����2�� #�#�"##�" �$5#� �$E#� O4U# � ^"� f"� o4u#� �~"���я�2xk[� 46�A��Q�P<��P�D�AՒ��HIuS}�zk[ ��� 2021-0�4-21�V � ;qb'_9_K_�]_o_�_�_�_�_�_ �L[T�Q18-02-27Y�_
oXo.o��T�8�:P�Qocouo�o�o�[N���W1�A�_�o�o�\��C���BX��; � `th&t92�@x�t�&t��'s���8�9�Jo� LM���hU��o����C<��D���-r:3�ErRqt�t�t�ht�2�@�t���.�RL�ڽh2��� ����5�r�%r�@-z��@92*pEz.�@�t�9�[��RK��hZ�;�z���r*pS!0's��ҟQ�������VJ�n�h�"a��N�`�r�r���ݍf�7���ʯUQ���n�-��G� �O_Z1 sM�_�q��� ������˿ݿ��_;��%�7�I�[�I`:�@c \χϙϫϽϫo�o���u��Bdp=�%p�d-p=��M�'�=� Ep=��M�UpM�]p�d(ߛ߉������� �v=������Z�t�;� �=��=��=҇�=� Q�=�Y��n������� ��ȍ��%p=�R�=�2 M�j�Q�c�u�5���J� \�������5�Mҹ�M� �������"4"�4� j|���������� ]���ާ�����L� �&�Z�|� ������/��@�/T/f/x/Ah�/ �/�/�/�/�/��9/&? 8?J?t҅P%r�P �P=p�2"��2��3��3]p�A�?�?�߿� ?OO�y7O �|;R Er�3R�P�P� P%��PY��O���? �O�O_ʍl?ZOlO~O �O4��_q��O�_�_�_ \?��oo�7oIo[o I[�o�o�o�_"_�` ���o�J�;��I_CFG 2{�: H
Cy�cle Time~�aBusyDw�Idlzr�t�mi8|�qU�pvv|qRead>�wDow8x�� �rqsCou�nt|q	Num Dqr�s�={��`�q��PROGWr|:D�0�u����������Ϗ�y �SD�T_ISOLC ; :� �@~�J23_DSP_?ENB  �>~#�INC }�|�e�A   ?OP�=���<#�
|�j�:�o u�������a��ȟ�OB�K�C,��uU��G�_GROUP 1�~�U�<� � �j�Cy.�П?"Dxd�m��`Q���� ��̯�����&�Dw���ڙG_IN_�AUTO�Q�#�P�OSRE���KA�NJI_MASK���t�KARELMON :(��by���(�:�L�@~�²O��V�X��xnŉ���CL_Ld��NUM0�����E�YLOGGINGĠ�?�v�U�F�LA�NGUAGE �:
��DEFAULT �6(LGXq�V��r��4�  �8�p��`'�g � ��`�ۏ�;���
��(UTg1:\\Ϧ� �� �����������!�8�E�W��(��#L�N_DISP ��M��x������OCgTOL���aDz@���f��GBOOK �)��z�qz�z�� 'Uy�k�}��� ��������5Ӱs����	-�t�*��/ُ�`�+�_BUFF {2�� A�Evꂒ�w� ����#,Y Pb���������/��ZDCS �V�Y�n���#�Dx^u�/�/�/�/6$I�O 2�B+ cp�/cp@���/?? *?>?N?`?r?�?�?�? �?�?�?�?OO&O8O�JO^OnO�O�O�O�%E_R_ITM��dD� �O_#_5_G_Y_k_}_ �_�_�_�_�_�_�_o�o1oCoUogo	��BS�EV�����FTYP���O�o�o�ovm΅�RST��4%SC�RN_FL 2�
�-@��g/gy�`����TP������b�NGNA�M,�`�
�2$UPS���GIp��U��B�_LOAD�G� % �%DR�OP��MAXU�ALRM�¢� ��U�
��H�_PRDM��� !���C���7�������P 2�7� �q�	�ol�W���{��� Ɵ���՟���D� /�h�S�������¯�� �ɯۯ��@�+�d� v�Y������������� ߿��<�N�1�r�]� ��yϋ��Ϸ������ &�	�J�5�n�Q�cߤ� ���߳�������"�� F�)�;�|�g����� ����������T� ?�x�c����������������DBGDEF� ��[!��_LDXDISA-���{�#MEMO_A�P'�E ? �
 $x(�����������FR�Q_CFG ���(A x'@�4E��<[$d%m�$:���^��*�/� **:����� _����+/"/4/a/ X/j/�/����/�@�/0�/�/�/�',(�/>? �$,?i?P?�?t?�?�? �?�?�?OOOAO(O�eOwO^O�O��ISCg 1� �� ��� �O��)�O��2__V_��O�B_MSTR ���myUSCD 1�o�N_�_J_�_ �_o�_4oo1ojoUo �oyo�o�o�o�o�o �o0T?xc� �������� >�)�N�t�_������� ����ˏ���:�%� ^�I���m�������ܟ ǟ ��$��H�3�l� W�i�����Ư���կ ����D�/�h�S���`w�����Կj_MK'���]Y�$MLoTARM&�-� 3" P�|X� METPUK �ǲ���YNDSP_ADCOLrż& }�CMNT�� ���FN���τ�F�STLI���ǁP ��^'�G�Y?�IԾ��POSCF�����PRPM��Y�S�T��1��[ 4Q#�
��ϱ���� �׿�������7��+� m�O�a�������������E�/��S�ING_CHK � ��$MODA�%��K���D�EV 	N
	�MC:��HSIZ�EKǰ��TAS�K %N
%$1�23456789�  2}�TRIGw 1��[ l�^9n�=Y�P��5��~�EM_INF 1���`)AT&�FV0E0�+)�E0V1&A�3&B1&D2&�S0&C1S0=>)ATZ+fH��:��bA�/�'//K/]/ �/5GYk�/ � ?7/$?6?�Z?? ~?�?w?�?g/y/�?�/ �/�/2O=?�/hO�?�O GOQ?�O}O�O�O
__ �?@_�?OO)O�_MO �_�O�_�_�Oo�_<o No5oro%_7_�o[_m_ _�o�_&]oJ o�;�����o ��o�o�o�oX�|� �����e֏������0���NITOR��G ?��   �	EXEC1T˳s�2y�3y�4y�Q5y�C {�7y�8y�9˳t��rޔx�ޔ ��ޔ��ޔ��ޔ��ޔ ��ޔ��ޔ̒ޔؒޓU2�2�2��2	�U2�2!�2-�29�U2E�2Q�3�3��3���R_GRP�_SV 1� � (7�5�(>����<�ȴ�0+&��=I?g�j���
_Dς���9�ION_DB���Ǳ  ���	��~���І�����v�W�&�N/   ?��?�����̢�-ud1�����υ�PL_NAME !�<��!Def�ault Per�sonality� (from FsD)����RR2��� 1�L6�L�A�<��� d:҉ϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻����������2��.�@�R�d�v�@��������<� ����0�B�T�f�x�����������޲�D����
���P J\n����� ���"4FX '9������ �//0/B/T/f/x/ �/�/k}�/�/�/? ?,?>?P?b?t?�?�?�?�?�?�?�> �H�6 H�b �H\���  �O1M�dC@PO bMFO�O�G@�=�|C��O�M�O�O C  �H__ _2_P_V_t_@�_�f��_�\��E�	`_�_o o�Q:�oA`�@oRodo�vn A�   �i�O�o�Lޱ�o�k�O �o'9$]H�: �R�� 1�4ɴ���R@ � �&�<��p @D��  �q?��s�q?���q�A��6E�z  �q���;��	l�r	 ��@� �0�ް!� ���p� � �� �F��J���K ��J˷��J� �J�4�JR�<g|v�f0O����@�S�@��;fA6A���A1UA��X{����=�N���f������T;f��X���ڀ��* � ��  �5'��>��p�H���?��?���{#�����ԏur`�f��q{��g�������i�V����(  ���������ʔt柉�	'�� � �I�� �  ���e��:�È(�ß�=���@���߶� <!��� � �  ��qz�˂�r�o�o����ү � '覵��@!�p@�a�@���@��@��C�C�"��"��B�pCz%����@�r��  ����n��������m;a;n�`@����D�u՟ҿ�� �����Q�c�E�U�ޔ�� :�W  }x�x?�ff�O�Ϙ�*� �P����⍁8�����>�A�x��q����0�P:��U�7�0�0���>����|���<2�!<�"7�<L��<�`N<D��<���,h��ߴ��s���s ҈`?fff�?��?&�аT@T����?�`?Uȩ?X�� ��L����t,��t8��w W�����ό�w��� ��������.��R���!�F�A���=����)���M����H�mN H[���G?� F��H ZE~i���� ��� �oAK ��������)�� �/��%/7/�j/U/�/y/�/�/��M��"�i��C�/?�/5? =�8��??F??j?���e��s��-M�BH"�E�.��?,�[2�Y0�X1�1@Iܔ=@�n�@��@�: @l��?�٧]�? ���%�n�������=�=D���0OB@��@��oA�&{C/� @�UXO��+J8��
H���>��=3H���_�O F��6�G��E��A5F�ĮE���O�@��f�G��E��+�E��EX���O�@>\�G�Z�E�M�F�lD�
�p�O�?E_ 0_i_T_�_x_�_�_�_ �_�_o�_/ooSo>o wobo�o�o�o�o�o�o �o=(:s^ ��������  �9�$�]�H���l��� ����ۏƏ���#�� G�2�W�}�h�����ş ���ԟ���
�C�.� g�R���v�������� Я	���-��Q�<�u��`�r���fB(hA43���h���൘��3�ϩп��!4� �{����!�0�+#(�:��jb�T�f�1E�䴛|�Ђˀ��Ϯ�����(���iP��P:�IVc߶�oߙ߄߽��ف����������9�$��"$<�N��r� �����v�H���&��e,�6�l�Z�|�����n)���������8F
  2 oH�6�&H�{�g\��&B�!�!� SB��0�0A� @�/ ��$�3���l^pUgy�T��$0� � ���� T�%
 ��//+/=/O/ a/s/�/�/�/�/�/�/�^J� ��$�����4�$MR_CABLE 2�$؟ � V�T*P��@n�?�0F1L�?0��0z Bz �C[0n�OM�`Bw���n��)��� D���G??Q6�  B�� TO�
�vr0����9���WD��2�h�?�7� �� C� ]9h4��r0��w�N~6���?��?�*\0�� [@CLW@j27�(Ԧn�:̉c�6E�/T3�O R˰O�O�O�O�O_�O �O"__*_�_�_`_�_ �_�_�_�_oAn�+��_Qocouol�?o�o��o�ol�*�o*�* 3OM ��%9��zH���%% 2345678901%�7u "RFqn�[@ j�n�n�
Lw��nnot segnt �jzsW,��TESTFE�CSALGRI�gDkʝd�t��q
�tG �P�n��"���'�9�K� 9U�D1:\main�tenances�.xmlS���  ���DEF�AULT2GR�P 2�	z  �pLn�  �%�1st mech�anical c�heckL}n��F6��>�G�H� $r���������n���controll�er��7��I�c�8�J�\�n���ϑ�M���n�"8��n�ȡϯH'�����*�<���Cٟn�����Y����ҿ�����ϒC�ge�.� batteryς�W�H	���ϖ��Ϻ���ϑSup�ply grea�sK���È�
�<���Hs�H�Z��l�~ߐ�ϑ �caCbl��߾�g�
7� ��0�B�T��ؑ+�����Q�����������`�$��@�hoo� ����������� +� O�a�s�)Zl ~�����'9  2DV�� �{����
// k@/R/�v/��/�/ �/�/�/1/?U/g/<? �/`?r?�?�?�?�/�? ?-?OQ?&O8OJO\O nO�?�O�?�?�OO�O �O_"_4_�OX_�O�O �_�O�_�_�_�_�_I_ om__To�_xo�o�o �o�oo�o3oEoWo >Pbt��o��o ���(�:�� �p��_����ʏ܏ � �O�$�6���Z��� ~�������Ɵ��9� K� �o�D�V�h�z��� ۟������5�
�� .�@�R���v�ůׯ�� ��п�����g�<� ����r����ϨϺ��� ��-��Q�c�8߇�\� n߀ߒߤ������)� ;���"�4�F�X�j�� �������������� �m���T���C���� ��������3�i� >��bt����� �/S(:Lp^p��	 T~ �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO�xO  �?�w  @� � �O�O�O��O__(_�*H_**  ���@zO|_�_�_b_p�_�_�_�_��! __�_Ko]ooo1o�o �o�ooo%o�o# 5oAk}��o�o Q���E�1�C� U����a�����ӏ�����	��e�w��
��$MR_HIST� 2��v�� �
 \�$ 23�45678901P����P�BR��9� ��������?�Q�c� �,�������t���ԯ ��ί;��_�q�(� ��L���˿��￦�� %�ܿI� �m��6ϣ��Z����ϐ���[�SK�CFMAP  ��y��Bʵ�����ON?REL  ��v��.�6��EXCFE�NB`�
,��y�F�NC��r�JOGO/VLIM`�dv��Ю�KEY`�����_PAN_����Ү�RUN����SFSPDTYP��<k��SIGN`�rԟT1MOT��o���_CE_GRP7 1��.�~� ��O��÷���a��� ���C�U��y�0��� ��f�������	��- ?&c���� t����M�q(�QZ_E�DIT]�(�Q�TC�OM_CFG 1��$������ }
�_ARC_}��`��T_MN_oMODE]���UAP_CPL/���NOCHECK� ?$� �� �/�/�/�/�/�/ �/??0?B?T?f?x?��?�?I�NO_WA�IT_L\���N�T��$�3����1_ERR��2�$�6ф�OEOWOiO�L�<юO�O�53 OC��#M| ��f�����A(C���$�8Ο,�C�#C3�ĳ�9<�� ?���_�O?�7NBPARAuMB�$���F�g�_yW8ѫ_�[ = ���_�_�S�_o(o o4o^opoLo�o�o�kxW��o�l}_n#�UM_RSPAC�E!��b�GQt�$?ODRDSP#_����OFFSET_�CAR�_/�vDI�S��sS_A3 A�RK]�OPEN_FILE�p_����cqPTION_�IO�����M_P�RG %3z%$�*A�S��sWO�p-����C쀄�\���  ;�?�r���g��	 ��ȴ�����4�dpR�G_DSBL  �n�.�J��sR�IENTTO_�f��C�>�-�A �r�UT_SIM_D��+ҋBdpVhpLCT ��=����O}��d\�_PEX�; ���RAT;' �d�����pUP S�m��pw����� �>�L��$PA�L�2��>`�_POS_CH�p��`�ZP�2��L6�LwA�W��� �oѯ�����+�=� O�a�s���������Ϳ�߿���'�9ϵ�2 ��h�zόϞϰ����� ����
��CW�4�F�X� j�|ߎߠ߲������� ��*
AAs'�}I5�4�Z�
BPG����� ��������&�8�J� \�n�����a�s����� ����"4FXj |��������� 0BTfx� ������///_�xW�Y/k-�� �c���/�+�/�/�'>-@>-�o?�/3?�'tP (7R?H?Z?l?�?�?�?��?&0w��?L�D(4	�`<?6OHOZOA:�o<�xO�O�O�O�`A�  �I!?�O �__�]?>_)_b_M_�__�_�_�_u����O��1������� ��$B@� �؄��P @oD�  a?�c��Q?<�a<�D� � Ez0c�:�;��	l&b	 ��@� �0PP_` ��
`� � �� ��b�PH0#�H��G�9�G�ģG�	{Gkf���GΈK/�o,�l�PC�1��`[��D	� D@ �D7g�n�d���  �5��>(p�`�4�(: �B4�Bp{{�!<���O��"��r'a�sW��Ao�Rҧpߐ��p(  ��p�����_$��U	'�� � B�I�� �  �<�E�F=���f�x�~��� <_`�� � ?� ��ف���8� b__�WN=��  'N�(��a�OpC�`��`[pB�`Cc5�G� ����@�i����m��A��G�MuAuN�@@<� �*b7e����4���X�C���������<�ȧ :�a�tx?�ff�/į֯h�C @��O�8<�<3�A�>�׶q"a�J�pn�Px���uanc<nd؃>������u�<2�!<"7��<L��<`N�<D��<��,0�o��c� c^���@?fff?�?y& �K�@T�2��?�`?Uȩ?X�B�:銒� 'd�Iev�g���Zd ���ϵ��������6� !�Z�l�Wߐߢ�y��� ����aσυ���D���HmN H[�ArG� F��M� ����������� ��(��%�^� _��� K�����+���g� *<N�cu� �����Β���I={C�O�s^?��}��,�?yç'c�'sqH�`�xp������:!@I��>}@n�@���@: @l���?٧]/ ���%�n��߱���=��=D��n/� ���@�oA�&�{C/� @��U�/ �+J8���
H��>���=3H��_��/ F�6�G���E�A5F�ĮE���/�� ��fG���E��+E���EX�?� >\��G�ZE�M��F�lD�
 `8?/�?n?�?�?�? �?�?�?O�?OIO4O mOXO�O|O�O�O�O�O �O_�O3__W_B_{_ f_x_�_�_�_�_�_�_ oo-oSo>owobo�o �o�o�o�o�o�o =(aL�p�� �����'��K� 6�H���l�����ɏ�� �؏��#��G�2�k� V���z�������韤"=(�!4�ퟦ�����֕3�ϩx� ��!4 �{:�<L��!�0+#f�x��Z�jb����1E�䴛|���������"��F�4���P޲Px���������@��׿¿��湿��π�A�,�Q�w�bϝ"$ zό��ϰ�����ߴ� ��@�.�d�R�ej�t���ߘߺ�������) ����.��R�@�v���  2 H�6f�&H�����\��&1B##B�  A� @'�����"�4�F�W���߁�������������$�R� � q�� ���%
 ��3EW i{���������* ���b����4�$P�ARAM_MEN�U ?����  �DEFPULSE��+	WAITT�MOUT�RC�V� SHE�LL_WRK.$�CUR_STYLv�OPT��N�PTB��C�R_DECSN� i�<,6/H/Z/�/~/�/ �/�/�/�/�/?? ?�2?[?VSSREL?_ID  ������j5USE_PR_OG %e%W?�?k3CCR�|2���m�7_HOST !e!�4O�:AT���?-C�?A/C|iO�;_TIME��|6�5VGDEB�UGz0ek3GINP_FLMSK�O��ITR�O�GPGA��@ �Lp� [CH��O�HTYPEbn�V?P?�_�_�_�_ �_�_�_oo?o:oLo ^o�o�o�o�o�o�o�o �o$6_Zl ~���������7��EWORD �?	e
 	�RS�@�PNS2��s�JO!��TEP@}�CO�L�3���3WL�0 U���	���5d�A�TRACECTL� 1���o� v�� �������&���DT Q嶾�S��D �� h�t��h� n�	 n�P$Pn� n��j��r��z���������n����l�l�	l���j��r��z�����������
l�l�l�l�k�}�������@şן�����`� :�L�^�p��������� ʯܯ&� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������ϰ
��.�@� T��T�|0V�T�T��T�T�T�T��T�T�T�T�(T�! V�T�T�� Z�l�~ߐߢ�쯮��� �8�J�\�n����\� ������������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ ���_�_
oo.o@oRo dovo�o�o�o�o�o�o �o*<N`r �������� �&�8�J�\�n����� ����ȏڏ����"� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����,�>�P�b� t���������ο�� ��_�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z������ ������
��.�@�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/�4/F/X)�$PGT�RACELEN � W!  ���V �l&_�UP ���e��!� �!� �l!_CFG ���%�#V!� ���$�$�/�'~ �*�  ��%�"DEFSPD ��,�U!~ �l IN~� TRL ��-��!8�%C1PE_C�ONFI� ��%O��!�$�)�l LID�#��-	~�9LLB 1�~7 ��$B�  B4�3�& �5JOE��/ << T!?�1KPO1OHOjO �O~O�O�O�O�O_�O��O_L_2_T_�_�Z B�_�_�_�_3O�_"o�o'oXo�9GRP �1��<W!@�  �[�V!A�?x�D P�DV�C2�� o�V d,D�i�i�1�0��0Wo)O�1�n#´(s
�kB+pRq�2.hR�V!>'oY>a�����~� =N�=R��3��0� i�T���x����Տ��x����  Dz0�9�V 
 �a��q��� ������ߟʟ��'� �$�]�H���l������)W!
V7.1�0beta1�$�ܠB(�A�?\)A�G��aޡ�>�������ޡA����f�fޢA�p��AaG��Q�Q@�(��`� ��K�]�o����#Apأ�r�0 ����Ϳ߿ڢU!��} ���v�$��H�2ϝ:�KNOW_M  ��%�&�4SV ���9��5 N�����f�9�$�6�Po��"�m�3Mvc����} ��	�%����T���P��$ߞ��פ�@ 1ߠ���(�wP�1+MRvcĥ�T~�D��u����OADB�ANFWD�ϡ3S�Tva1 1ś)��4�5�����& ��� �Q�D�V�h��� ������������
 O.@�dv������2�����V G�<%�w`3!3E��4bt����5������A6//,/>/��7[/m//�/��8�/�/�/��/��MA���d�3�'OVLD  �;�ߊ���PARNUM  �븆?�?��SCHS9 a5
�7�1�9��
EUPD�?�5uTO�%_CMP_��V0�����'��lDER_wCHKzE����0�ҎFwO�KRSg���Npa_MO���H_�O~�%_RES_G���;
8��oi_\_�_ �_�_�_�_�_�_o�_ /o"oSoFo9?+U6\F_xo+Ua�o�o�o -S��o�o�o-S  27-SZ Rqv-S � ���-S 0��<�-RV 1����ᾱ�@`z$�BT?HR_INRg�X1����dc�MASS6p� Z��MNo����MON_QUEUE ������@��U�$Nq@U�AN��ۈ�END��_��EXE ��6@BE����OPTIO���[��PROGR�AM %Պ%��.��?�TASK�_IU4g�OCFG� �Տ�?ɟ��D�ATA����@(�2��k�}����� ��^�ׯ�����ʯ�C�U�g�y�,�INFO���I���5�ҿ �����,�>�P�b� tφϘϪϼ�������@��(�:ߕ����I�� di���@DIT� ���߬���W�ERFLA�V���RGADJ Ή�/A�  ��?�@�w����� ��W�/�?���z��@'<@�9���%?h�0��dm�C�2�%糲+	H�l7�U�2�u?G�A ��t$���*��/�� **:���@������5,�'�����1��1W�9�Q����/�A� o�e�w����������� ��]G=O� s����5�� '�K]�� �/�����y/ #/5/c/Y/k/�/�/�/ �/�/�/Q?�/?;?1? C?�?g?y?�?�?�?)O �?�?O	OO�O?OQO OuO�O_�O�O�O�O �Om__)_W_M___�_ �_�_�_�_�_Eo�_o /o%o7o�o[omo�o�o�oN�	�<��*c Nt����Q�M����PREF ��%�����
��I�ORITY��܆�>��MPDSP������C�U������OD�UCT�������OG��_TG���钍ڂ�HIBI�T_DOA���TO�ENT 1Ӊ�� (!AF_I�NEm� �+�!�tcp+�S�!�udB�{�!iccmj�qXY��ԉ����)� 0��ߟ����ٟ� ��	�F�-�j�Q�c��� ��į��������$B�T�*����%����V����>rlD
�f��/	���������~��AG�,  ��o�D�V�h�(z��պ��Z뿺�������ϻ�i�EN�HANCE �u�s�A��d�P�7Մ~���������PORT_NUMn�������_C?ARTREP�Ĝ>�SKSTAm��oSLGS��ě��G�T�UnothingX�5�G��Y��{��TEMP �ڑ�e��e�_�a_seiban ���������"�� F�1�j�U���y����� ��������0@ fQ�u���� ���,P;t _������� //:/%/^/I/[/�/�/�/q�VERSI�L����  d?isablej�m�SAVE ۑ��	2670H7K55�(�/E?!@�0G?Y?|�}? 	�8w�$�o�;�?��e�?O"O4OFOTJ�<|?�Ot��5_�� 1�ě20�@r�e�O�O��g�pURGE�B掘�WFP�p�����W�3T�ѯ�W�RUP_DELA�Y ���&UR_?HOT %!vz��?߳_DUR_NORMAL�X���_�_�WSEMI�_�_;o�q_QSKIP�C�|��Cx�/�o�/�o�o�o �m}�o's�o!3E iW���w� ����/��S�A� c�������s�я���� ��ߏ�O�=�s��� ��]�����˟���>SRBTIF4T��RCVTMOU������/�DCR��C�^i ���aBJ�'B�[�yB��@�$��?(��)�����mH\�e���1��p����1R�oۯ�o �<2�!<"7��<L��<`N<D��<��9��O֯?�Q�@�u��� ������Ͽ�����)�;�o�RDIO_TYPE  �M�1�G�ED�T_C�FG ��KbB�HSE��Xa2�.� �ȸ��� ��.� �үD�/�h�S� �ϙ�(o���o��ӟ�� ���;�)�_�M��m� �ߴ�9�{�������� %��5�7�I����� ����a�������! E3i�����a� ]���A/ e���mG�� �/�+//O/qv/ �/G/�/C/�/�/�/�/ �/'??K?m/r?�/S? �?�?�?�?�?�?O�?�!OW?}?nO;���INOT 2�Y���_�G;� �O�K�+�<�OX�f�0 _[ 3O6_'OF_H_Z_�_~_ �_�_�_�_�_o�_2o o*ohoVo�ozo�o�o �o�o�o
�o.@& dR�v���� ����<�"�`�N����!�EFPOS1� 1�d�  x\O҉���O��� �+�ŏ׏�r�]��� 1���U�ޟy�۟��� 8�ӟ\�������-�?� y�گů����"���F� �C�|����;�Ŀ_� ��������B�-�f� ϊ�%Ϯ�Iϫ���� ߣ�,���P�b���� Iߪߕ���i��ߍ�� ���L���p���/� ����e�w�����6� ��Z���~��{���O� ��s����� 2���� ze�9�]� ���@�d� ��5G���/ �*/�N/�K/�// �/C/�/g/�/?�/�/ �/J?5?n?	?�?-?�? Q?�?�?�?O�?4O�? XOjOOOQO�O�O�O qO�O�O_�O_T_�O x__�_7_�_�_m__ �_oo>o�_bo�_�o�!o�o�oUc��2 1崏^opo�o(L Rop�/��e ����6���� /���{���O�؏s��� ����2�͏V��z�� ��9�K�]������� ��@�۟d���a���5� ��Y��}������ů ��`�K������C�̿ g�ɿϝ�&���J�� n�	��-�g��ϳ��� ��߫�4���1�j�� ��)߲�M���q߃ߕ� ��0��T���x��� 7����m������� >�������7������� W���{���:�� ^����ASe � �$�H�l i�=�a�� /���/h/S/�/ '/�/K/�/o/�/
?�/ .?�/R?�/v??#?5? o?�?�?�?�?O�?<O �?9OrOO�O1O�OUOx�O�o�d3 1��o �O�O�OU_@_y_O�_ 8_�_\_�_�_�_o�_ ?o�_co�_o"o\o�o �o�o|o�o)�o& _�o��B�f x��%��I��m� ���,���Ǐb�돆� ���3�Ώ���,��� x���L�՟p������� /�ʟS��w����6� H�Z���������=� دa���^���2���V� ߿z�Ϟ���¿��]� Hρ�ϥ�@���d��� �Ϛ�#߾�G���k�� �*�d��߰��߄�� ��1���.�g���&� ��J���n�����-� �Q���u����4��� ��j�������;�� ����4���T� x��7�[� �>Pb�� �!/�E/�i//f/ �/:/�/^/�/�/?�OT4 1�_�/�/ ?�?m?�?�/�?e?�? �?�?$O�?HO�?lOO �O+O=OOO�O�O�O_ �O2_�OV_�OS_�_'_ �_K_�_o_�_�_�_�_ �_Ro=ovoo�o5o�o Yo�o�o�o�o<�o `�oY��� y��&��#�\�� �����?�ȏc�u��� ��"��F��j���� )���ğ_�蟃���� 0�˟ݟ�)���u��� I�үm������,�ǯ P��t����3�E�W� ���ݿϱ�:�տ^� ��[ϔ�/ϸ�S���w�  ߛϭϿ���Z�E�~� ߢ�=���a����ߗ�  ��D���h���'� a�������
���.� ��+�d����#���G� ��k�}�����*N ��r�1��g����8?045 1�;?��1� �����/�/ Q/�u//�/4/�/X/ j/|/�/??;?�/_? �/�??�?�?T?�?x? O�?%O�?�?�?OO jO�O>O�ObO�O�O�O !_�OE_�Oi__�_(_ :_L_�_�_�_o�_/o �_So�_Po�o$o�oHo �olo�o�o�o�o�oO :s�2�V� ����9��]�� 
��V�����ۏv��� ��#��� �Y��}�� ��<�ş`�r������ 
�C�ޟg����&��� ��\�寀�	���-�ȯ گ�&���r���F�Ͽ j�󿎿�)�ĿM�� q�ϕ�0�B�Tώ��� ��߮�7���[���X� ��,ߵ�P���t��ߘ� �߼���W�B�{��� :���^����������A���e�K]6 1�h�$�^�����  �$��H��E~ �=�a���� �D/h�'� K���
/�./� R/��/K/�/�/�/ k/�/�/?�/?N?�/ r??�?1?�?U?g?y? �?O�?8O�?\O�?�O O}O�OQO�OuO�O�O "_�O�O�O_|_g_�_ ;_�___�_�_�_o�_ Bo�_foo�o%o7oIo �o�o�o�o,�oP �oM�!�E�i �����L�7�p� ���/���S���� ���6�яZ����� S�����؟s����� � ���V��z����9� ¯]�o�������@� ۯd�����#�����Y� �}�ϡ�*�ſ׿� #τ�oϨ�C���g��� ����&���J���n�	�x��x���7 1�� ?�Qߋ�	���-�3�Q� ��u��r��F���j� �����������q� \���0���T���x��� ��7��[�� ,>x����! �E�B{�: �^�����A/ ,/e/ /�/$/�/H/�/ �/~/?�/+?�/O?�/ �/?H?�?�?�?h?�? �?O�?OKO�?oO
O �O.O�OROdOvO�O_ �O5_�OY_�O}__z_ �_N_�_r_�_�_o�_ �_�_oyodo�o8o�o \o�o�o�o�o?�o c�o�"4F�� ���)��M��J� �����B�ˏf�� �����I�4�m���� ,���P���럆���� 3�ΟW����P��� ��կp��������� S��w����6�������8 1���l�~� ��6�!�Z�`�~�Ϣ� =ϟ���s��ϗ� ߻� D������=ߞ߉��� ]��߁�
���@��� d��߈�#��G�Y�k� �����*���N���r� �o���C���g����� ������nY� -�Q�u�� 4�X�|); u����/�B/ �?/x//�/7/�/[/ �//�/�/�/>?)?b? �/�?!?�?E?�?�?{? O�?(O�?LO�?�?O EO�O�O�OeO�O�O_ �O_H_�Ol__�_+_ �_O_a_s_�_o�_2o �_Vo�_zoowo�oKo �ooo�o�o�o�o�o va�5�Y� }���<��`�� ���1�C�}�ޏɏ� ��&���J��G�������?�ȟc��ҿ�M�ASK 1����0�>��XNO�  �=�C�MO�TE  _�  ���_CFG ������PL_RGANG������٦OWER ������SM_DRYPRG %���%��I��TAR�T �	�W�UME_PRO&�8�����_EXEC_E_NB  �����GSPD��ΰָ��TDB��R�M��I_AIR7PUR� ��m�\p��MT_�T������OBOT_I/SOLC]��l�̥�ȥ��NAME ������OB�_ORD_NUM� ?	�i��H755  ���@�R�d��PC_TIMEOUT�{ x�S232���1�`�� L�TEACH PENDAN�б�С���������Maintena�nce Cons�������"�ߒ�?No Use��� ��@�R�d�v������NPOf���С�����CH_Lf�����	�~��!UD1:1�z��R�VAIL!���������SPA�CE1 2�`�
��ХЩ�巓�ΦТ�m���<7 ���?�Y� Y���KlC�|�� �������%< �QrY`�d��� ���Y)/@/ �U/v/]/�/��� ���//7/-?�/Q? r?�?k?�/�/�/�/�/ �??3?)OJO	O_O�O gO�O�?�?�?�?�?O OAO7__[_|_�_e_ �O�O�O�O�O�__=_ 3oToou_�oqo�o�_ �_�_�_�oo)o/Mo e�]o�o�o�o �o�%G=�^�� ��{������� ��!�S�9����o����g������2��� ��ݏ����%�W� Z���:�������Ưǟ3ڟ����"�ԯF� x�{���[���ҿ����4����1�C��� g������|��������	�5�.�@�R�d� ߈ϺϽ�ߝ������)�*�6=�O�a�s� ��7������$���5��J�K�7^�p�� ���X�������E��� 5V-kl�8��� ������y�� f� VwN��G ;�� �ń�
� �   �//1/C/U/g/y/ ���-���/m�/ȁd0�/2?D?V? h?z?�?�?�/�/�.�: �?�;O??�?ZOlO ~O�O�O�O�?�?�?�? O_5_(O:O�Oz_�_ �_�_�_�_�O�O�O _�"_4o `� @Ȁme�/{oW__Y�a�UDo�o�o�_�j�o �o1CaI�� gq������ �Q�c���7�i������������Տ�ُ�\
��ol��A��*S�YSTEM*�V�9.10185 ���12/11/2�019 A ��� ��r�ӓSR_�T   � �$ĐENB_TY�P   $�RUNNER_A�XS� $HAND_LNGTH�`}�THICK���FLIPґ�`$�INTFEREN�CE��IF_CIH��I֑$�9��INDXD�ĐG1�POS   qW�N�`�ANG`��x�_JF��PR�M`� 	�RV�_DATAƑ � $��ETI�ME  ��$VA�LU����GRP�_   ���A  2 ��SCő	� �$ITP_�� $NUMڠsOUِ	�TOT��
�DSP!�JOG�LIM� $FINE_PCNT@��CO��$MA�X�TASK@�KEPT_MIR=�>]�PREMTq�}��APLD���_EX�������t�@��P�G��BRKHOL�D�!��I_� � ڲ@���P_M�ADE�w�BSO�C�MOTN�DUMMY163��SV_CODE_�OPM�SFSPD__OVRD��R��LDL�O�ORZ�T-PӐLE[�F!�[�6:�OV=�SF���ē�T�F��A�a�UF{RA��TOOL@��LCHDLYW�R�ECOVK��:�WaSs�:��=�ROM���I�_�ڐ @���S��NVERT.�OFS;�CǠD��FWDt���p��EgNAB��7�TR���`���E_FDO>��MB_CM���=B-�BL_Mi�]���Ҫ�2S�VSTAA�$UP�����G�׸�AM����а���%� �_M��A�A�M�A�1�T$CA�0�,�D�7�HB�K���L�IO?��[�IQ�$PPA O�{�`��s��s�1�?DVC_DB��F�����쑼��A���1���%���3��+�AT�IO� �h�K�U���/�/�P�ABF�T ֒E�G�Ԛ���E�:��_AUX�SUB�CPU�G�SIN!_7Ў���P�1�������FLA��ݑHW_C1���j������$ATR���$/UNIT�����ATTRI���G��CYCLC�NEC�A!�FLTR_�2_FIR�TAR?TUP_CN`Ӷ�oSIGNO�LPS��2�1�_SCTz�F�_��F_��t��FqSF����CHA���[���O��RSD�/���/�P��s�_T���PRO�|�p�E#MP�=��T����ܐ���'DIA�G�RAILAC4��p�M�LO�њ'�4�PS-�@� Xi�+�%�PR��SB�  �C�� �	$�FUNC����RINS_�TB���=�o�RA��`�7��a�E���WARq�8�BL'CUR�$A+	((DA��G(#%LD=�?�h�o#�2�to#TI��%��ܐ$CE_R�IA_SWA�AF���P^��#��%T�2\CK��CMO�I���DF_LEl�_�PD�"LM���FA�HRDYO,��E�RGt H� z����O 5MULSE�� ���0��$J�W�Jrǂ�FAN?_ALMLV�Î1�WRN�5HARD�אO�_O,� �2N�1STO�Ƶ_���AU��R�(���_SBR���5.�J����CMPIN�Fڐ��-De!8CREG@�NV0l�$��۱DAL_N��F9L����$M 2�Ȏ7%�ܐ�8�ECMj-�N0�Y���дG���SP$R�+$Y��Z����ۡ���� ���EaG!`
�?�
QAR��0�'�20�U3 ��A�XE$�ROB!�R�ED!�WR�߱_i]�SYܰDQᰋVS�WWRI�V���STR �)��f�E���Ġ&To�1�B��P1��V5c�OT�OHAĠ�ARY��b]�ΡR�FI���h�$LINK��!��3a$EXT)_�S1�%U6�[a�XYZ�2ej7sfO�FF9�2bZbNh`B���d�����cFI �g�A�47Ĩ9�_JL�¢@d�?ch��0�T�[8��US��B	qL2ArCL7 ��DUO�$V9pTUR�0X�#zu!ab(BX�P,�)wFL[`���@�P�p|e�Y30��G� 1ĠKF�M�'�3��s��8���a�ORQ.� ��x��s��m�� ��H��,�_A]�OVEd���Mh l��C~��C ~��B}��0{�B�|��� {�~��h� ��e�u� ����l�v�e�����C����.�ERK��	BtEЪ��E�A�ܐ�e� gN!K�N!AX�¢N!��� 4b��0��Z1��o�� `��r`���`��:p��qp��1�p��:0��:0 ��:0Ǚ:0י:0�:0 ��:0�:0�:0'�D��8�DEBU��$���3(�N�VbAB�NL�t�^�VA�� 
����+���7� 0�7�o7�a7�ra7� �a7�:q7�qq�$Fp�"\ۂ�cLAB�b)�����GRO: )r�<*�B_,��Tm� �`�0��*���1�AND�pt�:�+�_e=��1Y� *��A�Pm�0!|�- ^`NT�0���VELل��L~���SERVE��N�@ $�`�A]!��PO@ҹ ���`���@���!�@�  $�TREQ�r
 �tR
����"2�q I_ �	 l���[ERR�boI,��لNr�TOQلրLHPP���R�� G��%Ha���   �REP  �
 ,��#�=��݁RA�� 2	� d��s���� �@$r�� ̙���OC?!� � d�COUN�T�Q��FZN_C;FG	� 4��aF3T������ܣq ���o��@T��C �(�M��g2��0Ճ{����FA� ��&��XdP�����$SQ��G�dQPB��@�HEL}@Y�� 5pB_BA�S��RSR`F�"^SS��!M�1��M�U2p�3p�4p�5p��6p�7p�8��@�R�OO�p��V ]`NL��ALsAB��FN�A[CK�IN�Tg CU�0E0� 	_P�Udq�2ZOU��P��aH-�֨ �P��T�PFWD_KAR�w�iAf�RE��$0P8/`U!w�QUE`I  e�Up�r�0�1I�0��-�[`S��SF[aSE�M3��A�0A��S�TYSO� 	�D�I�}����!_�TMuCMANRQ�L[`END�t$�KEYSWITCaH^s.�HEUp�BEATM�PE�PLEv�����U�rF�sS3DO/_HOM� O�1 EFA�PR�a�vQ�P�EC�O01c��яOV_Mr� � IGOCMGt�A���v.�HK�A DXa$bG��U^ҹMP��W�WsFORCfCWcAR 2	P,�OMP  @��c�0U�SP3P1�&�@�$E3�&4����O� �L�"��aHUNLiO9 \�4ED�1�  �SNPXw_ASZ� 0�@�ADD��$S{IZfA$VA�~��MULTIP���.3� A�! � $H	/0��`�BRS}�ϱCrТ6F'RIFu��S� �)���0NFOODBU�P~��5�3�9�ƽAfIA�!$V�y�x�R��SN��@ � L0��TE�s8�:s�SGLZATAb�p&�o�sC᳍P[@STM�T�q�CPP�VBW<e�\DSHOW�Ev�7BAN�@TP�`�w@qs8��s8��r �V7��_G�� :p$PaCD �7���FB�!-PXSP� A U���VDP��w� �W�A00^� ZR� bW� bW� bW� �bW5`Y6`Y7`Y8*`Y9`YA`YB`Y�  bW��cV�@bWF`X7� $hlY(@$h�Y@@$h�YU1�Y1�Y1�Y1�YU1�Y1�Y1�Y1iU1i1"i2_Y2lYU2yY2�Y2�Y2�YU2�Y2�Y2�Y2�YU2�Y2�Y2�Y2i2i2"i3_Y�p�x�yY3�Y3�Y3�Y3��Y3�Y3�Y3�Y3��Y3�Y3�Y3i3�i3"i4_Y4lY4�yY4�Y4�Y4�Y4��Y4�Y4�Y4�Y4��Y4�Y4�Y4i4�i4"i5_Y5lY5�yY5�Y5�Y5�Y5��Y5�Y5�Y5�Y5��Y5�Y5�Y5i5�i5"i6_Y6lY6�yY6�Y6�Y6�Y6��Y6�Y6�Y6�Y6��Y6�Y6�Y6i6�i6"i7_Y7lY7�yY7�Y7�Y7�Y7��Y7�Y7�Y7�Y7��Y7�Y7�Y7i7�i7"d �VP�U� �߰e��
FQ�2�� x e#�R�@  ���M��R9� ��Q_�+�R����(�~ ��S�/�C�D�^�_U8�0i��"YSL���� � L5Bj��4A7�D����&RVALUj�% x1���=F��ID_L�3���HI��I�"$FI�LE_L!�i$������SA�� h	�M�E_BL�CK�Z�uAc�D_CPUs�M0s�A0u��$�6�-0YZ@FR � � PW�-����0��LA�A�S�������RUN_FLG���� ���@v�!���!���HF ���C���l1T2x_�LI�"  ���G_O�� P�_EDI�"D@T2��c�k�9��n���0�0 �TBC2LT �Q@ �(0�!c�FT���	TDC�A4z���aM�������TH�0"�!�#�$�R��0e ERVE�F�	�F�5A�� � � X -$q�L�EN�~�	q�) R1A� 2��W_?���i1q��2��MOk�5S�0 I. Z��0���q���DE�1�LACE,":�CC83Z¶_MA208>>TCVEfTXg
�|
8RP1Q�1QJA-U�M���J>JP�}�2��@0P�	0JKVK@�A.)A.5A#J�AlF2JJ:JJBAAL2h:hbdAAf5#� N1�P�XB G�L��_�An�0�����CF62�! `	�GROUP��vA�2$QN��C�3~�REQUIR1��0EBU�3m��$T 2 *!n�&8��50��" \� ��oAPPR  CLG��
$t�Ng(CLOD��w)S��)
��.u6# ���M �C 8� 2�$_MGA� �CLPN��(� R �'B{RK�)NOLD�&�@RTMOb�:
=�%Jb�4Pj  :�  B  �  �  6W57W5hAB�m��$� "���A��7)A�3PATH �7�1�3�1���3� / 9#\�PSCA�� 7lh"�!INp�UC����0@C:PUM9HY��?�� @A��L�[J��0[Jq0[@PAYL�OA7J2L�R'_AN��CL�ЦI�A�I�A�%R_F2�LSHR@��ALO��D~A�G=C�G=CACRL_��-E P)G�Dr�H��G�$H�"^NRFLEXj#Z�;BJ��% PT"����E�W���Jp�& :}��� �W��T��� ������F1�QEeYg������(�bE2DVh z����`x}t� �m`�x���QT�w^qXF�� �d�h%.�x1CU gktb����t�j�J�' ���`��	/���ATrf!� EL�`(�D�#(�J/ &* JE0C3TR)AmaTN��@��'HAND_VB�G�jQ���4( $��pF2�&���S�W�#�&)� $$M�@�)!��!�@1�#p��E2�A�� �@�&��<��-A�,��
�*A;A;G��+�Ъ�*D;D;P�0G��ݩST�'�9�N8DY�e �&(� O��@r��G�Q�G�A�G �t`�5P_5h5�q5z5�5�5�5�2RD�R�4* ��T�2� �a㵙!�AS�YMEZ� F)K� L�A$O_B�X5@ HD2=4ĸ�ROdOvO�O�CJ�LR0�J�����I.d_VI��ؙ#!�V_UN���6�W��AJN�|�N��L R�U_ԃ�]� $YR0�3_E_���[TcS � ���HR���a+���}P]"DI0�#O#����,) g�V�I9�AV1S P�s`^�^�v`���`� - � ɑME�a��y���`�T�PT��Հ�0����V ��������T��� $D�UMMY1q1$7PS_p`RF2`���$���PFLA��YP���$GLB_T��1����]!�0�`q�}�. �XT '�1ST��* SBR�0M21�_V&"T$SV_�ER�@O��w��C)LK�w�A�`OS� ��GL�EW�/ �4���$Y��ZB��W���AœAz�9BΥ0��U��0� �pN���$�GI��}$�� �������1 L����}$F��E^NEAR�`NwcyFd	�`TANCwb���JOG&`H0 �2�P$JOIN�T�"�����MSE]T�3  EJ�a�S�� 1��_4� n`U�a�?�* LOCK_�FO�@Б�BGL�Vt�GLTES�T_XMj �EM�P� &"2I�� c$U�P��9`20* ���X1#̐� X/�y�CE�&y $�KAR$qM%�TP�DRA���VE�C`�� IUX2�]HE TOOL�9c�V8dRE�I�S3�U�6z1m`ASCH� / 3�O@ԩ���3g�% SI�Z"  @$RAIL_BOXE����ROBO)?����HOWWAR�VQH!��!ROLM �n%ԁ$"�6 a`n�0O_F�!��HTML5�)A�Ͳ��!�15��R�O�R6�"1`�ئ ���OU�7 	d��T/`�J�$�� _$PIP*N�p��6"!`X� �PCORDED� 
@� &a XT*0) � ��O`� 8 D 0�OB|�N�� �7�v1��/�v2��P�SYSv1ADRO� ���TCH� 9 M,�pEN	�QA�_�4݁�R��V�WVA|�: �� ����PRE�V_RT��$E�DIT(FVSHW�R�c�G@�b����D��O�^DW�$HEAD����x@���0CKE����C�PSPD�FJMP��0L��R�`;�Q;~0{Q�6I3SO��C��NE�P���T'ICK9c��M�Q�p��EHNY�< @p�0�AᅗA_GP&V�-&�PSTY�2!L�OK�N�B"R�P=� t 
#@G�5%�$A=c�SE�!$D�9`���M��9P&�&VSQU�,e<��TERC��ʱz�S�>  �o���p��q�``O����{`IZ����PR\0�Db�A�0PU;�Te_DO�i�0XS� K�A�XIs`�#]UR ��cP�O P�6���Y_��2ET�bP��0	�rPF	�sPA,����9'[�) ��SR��?l�P�!���/u�Ay �/u*�/s8�/sH�uu j�uuz�uu���u�}����u�|���yC
��}C��}�ϕϧϹĠ�SS}C3� @ h��cDS4P���SPJ�&��ATx� �UaP��B��ADDRESz�B3@SHIF�^O_2CHO��1�IR���TUR�I��� A�"CUS�TO�dP�V�I�>�B�2��8c�
.2
6�V1daN~�C \a�8�rPC�a�P��C��b�b�R�6���TXS�CREEx2D��QTINA��# Ӕ��#Q_��ٰE T�A��8b�1��n�� ��a�2�b�/@RROS�~ �0�@�o�� ;UE�DF ���1r
�S��1RSMP�wgUe0�P抡�S_��=Ú���ȧ=��aC���� 2-EΐUEմGD��\�D`GMT��Lp���a~�O��@BB�L_ W��~�H ��rPJ�O��V�L�E�a�N �`�RI;GHj�BRD��ہOCKGR����Tf0|����WIDTH#�T@�b)!��T��UI� EY��}�I�
2� m VR6 @aB�ACKTQ�Ũ���FOS1�LAB�_q?(��I �$URT!E���ް��}H@� J 8��B~ _wA�h�R�� �s(��R�O�~�%KP����Uv���9Ry!LUM�Øf�ՀERV!1��ްP�h �L���`GE`I�O�`l2�@LP��bE�Pf�)%�v�3�P��3�  2�50�60�70�8��R��?`h ����� !�S�P�KݱUSR��M <a���U(�sFO�PRI�a�m  ���TRIP�2!m�UNDO
;�N �P �ye`!�xeS�P�`�P O�c���CaG PT0� T��^�OS��s�AR�`F�J��Z�P��@������6T� OU�Z�Q���ã�5UJ�OFF([�R_�z��O)� 1P���;�Q��GU�1P�:��"V�Q�`��SUqB6R��i�SRT���tSR}� #cOR� ��RAU(p��Tȼ��7��_&@�DT 9|1p�8OWNM��4$SRCQ�Ҡ�P�D(&rMPFI8MT|��`ESPPab ����eA��������A@
�U `��WO�[p�4a�PCOP&��$�`O�_- bX�1�WA3@CF �� Z��p@l"�+� V�SHA�DOW�`��_UNSCA��ʴ�DGD!�1EGAC�8�� CWp`
�W� ,"w1�S$NER�c�Q�#+�C0cDRI5V6f�a_V/P���@m D��MY_UBY��kyV��UR���P�eA�h "P�_MT"LZkBMv]�$�@DEY�3cEX7�^��MU�@1X]�V$��US���`�_R�����
�R����G�pPACIN�A�PRG�$�"�`�"��"ң�RE}遚�c�H�"@XS �� G�P��H� �0IR��@Y���?�ӱ��	�qaRmEb#SW� _A�!�e�W#B`O��ہA(�^3/rE��UeP�d���IHKjRZ��v:�P&q[0%��3EAP�7� j�^5��IMRCV
�[ U��OvPMj�C���	�2��#�2REF 6�F�6�1M0���c50 ���:FAJFAKhE�6��?_ �:�H�;�pS���N'�aYUI�\ �GR�ӵ`�м�POU4W�"VkO W 5U�2��a$Ԑ��C`,�Y���U�2Q{�ՀULj��Z_ CO~��[H EPNTZ�Th�U ���V�ђSQPL��U�#�U���W���V�IA_���] ���`HD����$J�O��6��$ZO_UPL�W�Z|p�W!e�QPSp�0�_L=I��$EPEQ��k�a�QǑ΁��΀
��P]m�^� 0贃�a� ��CACHLO:A�d�aI оi��� 1CI`MI�FHa�eT�p�f�K�$HOj��`C'OMM���Ot�w�WӲ�S&�T7 V�P�"$Pmr_SIZwtZ� rx!asw�v��MP�zFAI!`5G�4�`AD�y��MRET�r|wGP���> & �ASYN�BUF�VRTD��%�|q��OL�Di_��A�W��PC���TU7#�`Q{0	�EwCCU�(VEM� x�e���gVIRC�q�9�!���%�_DEL�A�#&Q���AG:5�RK!XYZ̠��K!W1��8A��򱦀TN8"IM߁8���|���eGRABB��QYb"�f�_����LAS��r1�a_GE�e`u�&��;����T/S&N` ���%I����"ņ�BGf�V5��PK� ǆ�aWKGI��N#�`2F�@��`�qq�a+�aS��p�fN:�@�VLEX��b�����;��Nq��I? �-|�P� |�.$�3����- �"c��b�t�ĸ���a�ORD����1��w�RN�d $.MPTIT� �C�8�F�VSF����e  -�[�QK UmR�6SM!�f+���ADJ�N%�PZ�D>�g DƨBaA�L+`�p�AbPER�Is`��MSG_Q9�$}q�u���b��h+�"�g�J`�3p/�XVR#�in�b��T_OVRi��/ZABC��j�";s/@
�QZ]�#�kL+�=$L�-Bk_ZMPCF��lH���A����LNK�c�
 ����m� $,q�0��CWMCM� C�C����DP_A+A$J����Dbq�� �h �h ����
D��F�UX���UXE ]!f��	�]��]�o�p��oё���FTFsQ�Ӿ�r1	�Zb�gn {�}� ����YJ`D�� o�Y�R�pU�$H�EIGH�#"�?(�MP�.A�����Dp� � EX�$B�QPx �SHIF,�s��RVI`F��/B|�0�C`�dTF @{"�������WuD��_TRACE��V�A}��SPHER� q ,MP�)�;��$R�!p��� ���F���� 6�S|��F��  S�Px�2p������s���r�����	��U��C�ADC��8{l6�R  d� � ZD �Qx0C���a�l�l0�| ��6�V��@ 2|F���� D��P�����	�	F�, :$ZH~l�� ����� //D/ 2/h/V/x/�/�/�/�/ �/�/
?�/??.?d? R?�?v?�?�?�?�?�? O�?*OONO<OrO`O �O�O�O�O�O�O�O_ _8_&_H_n_\_�_�_ �_�_�_�_�_�_�_4o "oXoFo|ojo�o�o�o��o�o�oF��$SA�F_DO_PULSC�G��k�$qp�ď�|k���5qR ���`��XP������
����P��s��tq � �������*��<�N�`�r�����.�  ��2��tq��d��ȁ�rs�� @������*��܉�� � 6��/_ @J�TY J����������T D��������)� ;�M�_�q����������˯ݯ��~�����M�_�$��sNR�;��f����p���
�t��Di��q��  � ����R�q |ulq���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w������S��G����� ��0�B�T�f�x��� ��������������@"4FK��b0E� ҳD�ܽ����� �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?��?�?�? �?�?�?�?	OO-O�� QOcOuO�O�O�O�O�O �OLz��!_3_E_ W_i_{_�_�_�_�_�_ �_�Yoo,o>oPobo to�o�o�o�o�o�o�o (:L^p��������ø� �Ǔ�6�H�Z�l�~� ������Ə؏����  �2�D�V�d�#�m�\����������i�	12345�678ݲh!B�!ܺTz1!���
��.�@�R� d�v�������"�ïկ �����/�A�S�e� w���������ѿ��� ���)�;�M�_�qσ� �ϧϹ��������� %�7����m�ߑߣ� �����������!�3� E�W�i�{��L߱��� ��������/�A�S� e�w������������� ��+=Oas ������� '9��]o�� ������/#/ 5/G/Y/k/}/�/N�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�/	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_BS��]_�o_�?�_�_�_Ԛ�Cz  Bp�z �  ��2��� } �X
g_�  	��R2U_ <oNo`oro�l��\�+o�o�o�o�o" 4FXj|��� �������oB� T�f�x���������ҏ �����,�>�P�b� t����������Qa:�R<Ք ˕a?  ������#a#at  ��P#�;���`�$�SCR_GRP �1�*P��3 � ��R� �U	 _����� �����Qԑ�U������pٯǯ ��]�`6��C�,����m���C����lLR �Mate 200�iD 56789�0!`LRM|� 	LR2D ��~�
1234���Ц�d��hbճ ���}�ݣ}��cԑ����ѡ�	j4�F��X�j�|τ���#H���Ē�}��πį������̦<��1���A���e��WV��Vh�`,R��  [W��B��Pư�Ȯ��Ԫ�A�P��  1@�0�ժ�@�����# ?4���H�P'���ڪ�F@ F�`Q�Y�P�}�h��� �����������ʩ�р���J�5�G�Y�k�B�y���������� ��=(aL�p ��o�
'�����WA`�.4�@4�O>�7�4̧@��0n�PQ�����ݣT_��A���$����aĲ�1A 
/1/C/Q*!f(Hr/�/S/�P�#
b �/�/�/� ?�/$?,4�]�ECLVL  �1����>1�L_DEFAUL�TF4������0Z3HOTS�TRf=�z2MIP_OWERFE0�Uzr5�4WFDOg6� r5=2RVEN�T 1M1M1�3� L!DUM_�EIP,?H�j!AF_INEf0<+O3D!FTOZN�!O~O!�ϣO ��mO�O!RPC�_MAIN�O�H�8�O_�CVIS�O�Iy�_b_!TPUP�PUY_IdQ_�_!�
PMON_PR'OXY�_Fe�_�_�uR�_Mf�_Fo!RDM_SRVGorIg5o�o!R��d�oHh�o�o!
�@�MoLi�o*!?RLSYNC+Qy�8v!RO�S O�|�4e�!�
CEwPMTCO�M�Fk��!	��rCONS�Gl��Z�!�rWAS�RCaoFmI���!��rUSB��Hn ���O�Uc���?� d�+���O���s�П87�RVICE_KL� ?%�; (%�SVCPRG1�ן�	�2�$��3�G�L��4o�t��5������6��į�7@�����/�*�97�<���od����� �9����a�ܿ��� ����,��ٯT�� �|��)����Q��� 6�z���6����6�ʿ D�6��l�6�ϔ�6� Bϼ�6�j���6���� 6���4�6���\�^�
� ܟ���������.� �����8�#�\�G��� k��������������� "F1X|g� �����	 B-fQ�u�� ���/�,//P/ ;/t/�/q/�/�/�/�/ �/�/??(?L?7?p?��_DEV ��9�UT1:�|?�0GRP 2
��5���bx 	�� 
 ,�0 x?�?�2�?OO@O'O 9OvO]O�O�O�O�O�O �O�O_*__N_5_r_ �_�?�___�_�_�_o �_&o8oo\oCo�ogo yo�o�o�o�o�o�o 4�_)j!�u� �������B� )�f�x�_��������� ����M�,��P�7� t�[�m�����Ο��� ��(��L�^�E��� i������ܯ�� �� ��6��Z�l�S���w� �������ѿ���2� D�+�hϿ�]Ϟ�U��� ����������@�R� 9�v�]ߚ߬ߓ��߷� ������*��N�`�G� ��k��������� ��&�8��\�C����� y���������C��� 4F-jQ��� �����B )fx_����� ���/,//P/7/ t/�/m/�/�/�/�/�/�?�/(??!?^?e3d �e6	L?�?�?�?`�?�?�?OK%�O<5O<C���NA�1 NE^OlGVO�OzO�O�O �O�I"O_JI�O4_"_ X_F_h_j_|_�_�O�_ _�_o�_0ooToBo do�_�_�o�_�o�o�o �o,P�ow�o @�<����� (�jO�����p��� ����܏ʏ �B�'�f� ��Z�H�~�l������� ؟���>�ȟ2� �V� D�z�h�����ůׯ�� ������.��R�@�v� ����ܯf�п���� ��*��Nϐ�uϴ�>� �ϖ��Ϻ�������&� h�Mߌ�߀�nߤߒ� �߶���.�T�%�d��� X�F�|�j������ ��*�����.�T�B� x�f������������ ��*P>t�� ���d���� &L�s�<� �����/T9/ K//$/�l/�/�/�/ �/�/,/?P/�/D?2? T?V?h?�?�?�??�? (?�?O
O@O.OPORO dO�O�?�O O�O�O�O __<_*_L_�O�O�_ �Or_�_�_�_�_oo 8oz__o�_(o�o$o�o �o�o�o�oRo7vo  jX�|��� �*�N�B�0�f� T���x�������&� ����>�,�b�P��� ȏ����v���r���� �:�(�^�����ğN� ����ȯʯܯ� �6� x�]���&���~����� Ŀƿؿ�P�5�t��� h�Vό�zϰϞ���� <��L���@�.�d�R� ��v߬�����ߜ�� ���<�*�`�N���� ����t��������� 8�&�\������L��� ����������4v� [��$�|��� ��<!3�� T�x���� 8�,//</>/P/�/ t/�/��//�/?�/ (??8?:?L?�?�/�? �/r?�?�? O�?$OO 4O�?�?�O�?ZO�O�O �O�O�O�O _bOG_�O _z__�_�_�_�_�_ �_:_o^_�_Ro@ovo do�o�o�o�oo�o6o �o*N<r`� ��o����&� �J�8�n������^� ��Z�ȏ���"��F� ��m���6��������� ğ����`�E���� x�f������������� 8��\��P�>�t�b� ��������$���4�ο (��L�:�p�^ϔ�ֿ �������π���$�� H�6�l߮ϓ���\��� �������� ��D�� k��4�������� �����^�C����v� d�����������$�	 ������<r`� ����� � $&8n\��� ����/� /"/ 4/j/��/�Z/�/�/ �/�/?�/?r/�/i? �/B?�?�?�?�?�?�? OJ?/On?�?bO�?rO �O�O�O�O�O"O_FO �O:_(_^_L_n_�_�_ �_�O�__�_o o6o $oZoHojo�o�_�o�_ �o�o�o�o2 V �o}�FhB�� �
��.�pU��� ��v��������Џ� H�-�l���`�N���r� ������ޟ ��D�Ο 8�&�\�J���n���� �ݯ������4�"� X�F�|������l�ֿ h�����0��Tϖ� {Ϻ�DϮϜ������� ���,�n�Sߒ�߆� tߪߘ��߼����F� +�j���^�L��p�� ������������� $�Z�H�~�l������� ������� V Dz�����j�� ��
R�y �B������ /Z�Q/�*/�/r/ �/�/�/�/�/2/?V/ �/J?�/Z?�?n?�?�? �?
?�?.?�?"OOFO 4OVO|OjO�O�?�OO �O�O�O__B_0_R_ x_�O�_�Oh_�_�_�_ �_oo>o�_eowo.o Po*o�o�o�o�o�o Xo=|op^�� ����0�T� H�6�l�Z�|�~���Ə ��,��� ��D�2� h�V�x�Ώ�ş��� ����
�@�.�d��� ��ʟT���P�ί��� ��<�~�c���,��� ������ʿ�޿�V� ;�z��n�\ϒπ϶� ������.��R���F� 4�j�Xߎ�|߲����� �ߢ��ߞ��B�0�f� T���߱���z����� �����>�,�b���� ��R������������� :|�a��*�� �����Bh9 xlZ�~�� ��>�2/�B/ h/V/�/z/�/��// �/
?�/.??>?d?R? �?�/�?�/x?�?�?O �?*OO:O`O�?�O�? PO�O�O�O�O_�O&_ hOM____8__�_�_ �_�_�_�_@_%od_nQ��$SERV_M�AIL  nU�d`�JhOUTPU}TYhoP}@NdRV 2�V;  g` (�Q4o<�oNdSAVEzlhi�TOP10 2>�i d j_  2DVhz��� ����
��.�@� R�d�v���������Џ ����*�<�N�`� r���������̟ޟ�0���U�eYP�oKc�FZN_CFG ;�Ugc�d��a�eT�GRP 2�^��a ,B �  A��nQD;�� B���  B�4�cRB21��fHELLW��U�f�`�ou���%RSR��)� b�M���q�����ο�� ˿��(��L�7�p���ϔ��  ��a%�����Ϣ������oP��������Ǫ�2oPd����ɦ�HK 1׫ ߈߃ߕߧ����� ������%�7�`�[�m�������ìOMM ׯ�Ȣ�FTOV_ENB�Yd�a�iHOW_R�EG_UI7�LbIMIOFWDL�����l�WAIT�4���v���t`X�ܡd��TIMX������VAX`��l�_�UNIT3��iL]CQ�TRYX��e�N`MON_AL�IAS ?e��`heo���� �
t��#�G Yk}�:��� ���/1/C/U/g/ /�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_OqOO�O�O �O�OvO�O__%_7_ �O[_m__�_�_N_�_ �_�_�_o�_3oEoWo ioozo�o�o�o�o�o �o/A�oew ���X���� ��=�O�a�s���� ����͏ߏ����'� 9�K���o��������� b�۟������"�G� Y�k�}�(�����ůׯ 鯔���1�C�U� � y���������l���� 	��ƿ?�Q�c�uχ� 2ϫϽ������Ϟ�� )�;�M�_�
߃ߕߧ� ��d�������%��� I�[�m���<���� �������!�3�E�W� i����������n��� ��/��Sew�����$SMO�N_DEFPRO�G &����� &�*SYSTEM*ܢ� 	�RECALL ?}�	� ( �}0c�opy mdb:�*.* virt�:\tmpbac�k\=>192.�168.@07:?15032 IZ�l~�}5!fr�s:orderf�il.dat-e�mp;2544 �W��/}-�*.d���a/s/�/��
xyzrate 61 ,/>/P/�/�/?��'�/� @�/�/c?u?�?�1!�:prog_1.tp�/�S?�?�?O�8��5�YOkO}O�/!<O4:RO�O��O_�3x!D:\ �O+P�O�0�Of_x_�_
�4!Ua)_;_�9�_ �_�_O"O4O�_�_io {oo�O;o�OVo�o�o� }6!o�?1052 �oi{.!/;MxP��� �/�/��_�q����!?J{A�S������9!3o��ԁZ�l� ~�� ;�J{R�������T!�3?1.1?5:8892�`؟i�{��,�;�M�O� ����)���ͯ^�p������J�?�Q�����ϙtpd�isc 0��2 ���Ͽ`�rτϗt�pconn 0 �*�<�N������� 11 �Ͼ���a�s�8�ߘ{�1ick�?=��P�������drop�߿���b�t�<�2+�P�������1�Ͻ���`�r����� ��;�M������'� ����\n�����7 I���#�� �j|��3EW��/}7!�3�� ;�Z/l/~/>/�� R/�/�/?�2!_�_ G��/e?w?�?Z�_:? L6V?�?�?O/0/�/ T?eOwO�O�/7O�/RO��O�O_��$SN�PX_ASG 2����,Q�� P 0 �'%R[1c]@�_WY?��%W_�_f_�_�_�_�_ �_�_o�_7oo,omo Powo�o�o�o�o�o�o �o3W:L� p�������  �'�S�6�w�Z�l��� �����Ə����=�  �G�s�V���z���͟ ��ן��'�
��]� @�g���v�������� Я��#��G�*�<�}� `�������׿��̿� ��C�&�g�J�\ϝ� �ϧ��϶�������-� �7�c�F߇�j�|߽� ������������M� 0�W��f������ �������7��,�m� P�w������������� ��3W:L� p������  'S6wZl� ����/��=/  /G/s/V/�/z/�/�/ �/�/?�/'?
??]? @?g?�?v?�?�?�?�?��?�?#ODTPAR�AM ,U�6Q �	�'JP�'D�@'H~D��-PPOFT_K�B_CFG  �fC2USOPIN_�SIM  ,[�sF�O�O�Ov@=@RV�NORDY_DO�  }E�ERQSTP_DSB�N�sBU_aX=@SR ��I � &ȃE�_�\�T�CTO�P_ON_ERR�_;B�QPTN ��E�P�C��RRING_PR�M�_0RVCNT_�GP 2�E�A�@x 	Q_Poh@>o�wobo�olWVD%`ROP 1LI�@�a xI�g�o�o�oE BTfx���� �����,�>�P� b�t�������яΏ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�]�Z�l�~��� ����Ưد���#� � 2�D�V�h�z������� ¿����
��.�@� R�d�vψϯϬϾ��� ������*�<�N�u� r߄ߖߨߺ������� ��;�8�J�\�n�� ������������ "�4�F�X�j�|����� ����������0 BTf����� ���,SP�bt����bPRG_COUNT�Fs��R�ENBo��M��D/_UP�D 1{[T  
�gBR/d/v/�/ �/�/�/�/�/�/?/? *?<?N?w?r?�?�?�? �?�?�?OOO&OOO JO\OnO�O�O�O�O�O �O�O�O'_"_4_F_o_ j_|_�_�_�_�_�_�_ �_ooGoBoTofo�o �o�o�o�o�o�o�o ,>gbt�� �������?� :�L�^���������Ϗ ʏ܏���$�6�_� Z�l�~�������Ɵ������_INFO� 1@%& H�	 �c�N����r�?�2@B?�z=��t���"�DA�/�?������µ�B�QQ���=�@ @G� A�i��>�| >���� �D�b�����B��B�3�~ՠS�B�����²�B����j�r7菟5B��/��Y?SDEBUG�A ���d))Q�SP_�PASS�B?~c�LOG =�]J!  �����  �%!�UD1:\��#���_MPC��@%�#ϒ@!̱A� @!�SAV ���y�ظ�вC�׸SV��TEM_TIM�E 1��K � 0  ����C�CȀ�	��MEMBK  @%�%!����%�7�G�wX|& � @G���iߎߞ�b��߲����^� y�@ ����*�<�v�T�f�`x������ ��� ����
��.�@�R�d�v��e���������� ��(:L^p ������� ��SK�����@hRdX�� "�Q2sߣ�P�� �� �������%/7/I/[/O�u$� �u/���@�/�/�/���/�À?@'?9?K?]?o?�$s?�?���?�4^�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__�)�T1SVGUNwSPDy� 'c���4P2MODE_?LIM ��g�20T2=P]Q��/U�ASK_OPTI�ONX��g��Q_�DIr�ENB  ���c��QBC2_?GRP 2#c�0���_�"� C�c(\�BCCFG !��[~� o"Ekem`eo���o�o�o�o �o�o�o?*c N`������ ���;�&�_�J��� n�����ˏݏ��ɋ�� ɏ*�<����r�]��� ����H�ڟԯ��� ��,��P�>�t�b��� ����ί������ :�(�J�p�^������� ��ܿʿ�� �6�� �J�\�zόϞ���� ���������.�@�� d�R߈�v߬ߚ߼߾� �����*��N�<�r� `����������� ��$�&�8�n�\��� HϪ���������|�" 2XF|��n ����� 0fT�x��� ��/�,//P/>/ t/b/�/�/�/�/�/�/ ��
??:?L?^?�/�? p?�?�?�?�?�? O�? $OOHO6OlOZO|O~O �O�O�O�O�O_�O2_  _B_h_V_�_z_�_�_ �_�_�_�_�_.ooRo ?jo|o�o�o�o<o�o �o�o<N`. �r������ �&��J�8�n�\��� ����ȏ���ڏ��� 4�"�D�F�X���|��� hoʟܟ������B� 0�R�x�f��������� �ү���,��<�>� P���t�����ο��� ��(��L�:�p�^� �ςϤϦϸ������ ȟ*�<�Z�l�~��Ϣ� �߲�������� ��� D�2�h�V��z��� ������
���.��R� @�b���v��������� ����N<r (ߊ����\��8&\Fz��$TBCSG_G�RP 2"F�  �z� 
 ?�   ��������@5//Y/k+~�$��d@ ��!?>z	 HBLk(z��&j$B$  C�`��/�(�/�/Cz�/�(=A�k(333?&ff?��i%�A��/m?80 k(c�͎6S5�0DHp?�=@�H0j%K1�5j$�1D"N!�?�?�?�? ;OJ�(I&�(nE�OLO ^O�O�O�O�O�O_ [��H:Q	V3.�00�	lr2d S	*\PTTy�k_*_ �Q�I 8�Pt]�_  �_�_,�[~J2�%�=Q�o�UCFG '�F� �"j��Lb�ROlwl�wo�o�jO�o�o�o �o�o=(aL ^������� ��9�$�]�H���l� ����ɏ��Ə���#� �G�Y��� d�v��� 2�����˟�ܟ� � 9�$�]�o�����N��� ��ۯƯ��zf6� BF�H�Z���~����� ؿƿ����2� �V� D�z�hϞόϮϰ��� �����
�@�.�d�R� tߚ߈߾߬����ߴ ����>�`�N��r� ����������&� ��6�8�J���n����� ����������"2 4F|j���� ���B0f T�x����� /�,//P/>/`/�/ 0�/�/�/l/�/�/? ??L?:?p?^?�?�? �?�?�?�?�?O O"O HOZOlO&O|O�O�O�O �O�O�O_�O_ _2_ h_V_�_z_�_�_�_�_ �_
o�_.ooRo@ovo do�o�o�o�o�o�o�o *�/BT� �������� 8�J�\��l������� ��ڏ����ʏ4�"� X�F�h���|�����֟ ğ���
���T�B� x�f���������Я�� ���>�,�b�P�r� t�����6Կ����� (��8�^�Lς�pϦ� �������� ߾�$�� H�6�X�~ߐߢ�\�n� �������� ��D�2� T�z�h�������� ������
�@�.�d�R� ��v����������� ��*N`
�x� �F���� $J8n��Pb ����/"/4/F/  /j/X/z/|/�/�/�/ �/�/?�/0??@?f? T?�?x?�?�?�?�?�? �?�?,OOPO>OtObO �O�O�O�O�O�Ol� _._�O_L_^_�_�_ �_�_�_�_ oo$o6o �_ZoHojolo~o�o�o �o�o�o�o2 V Dfhz���� ���
�,�R�@�v� d���������ΏЏ� ��<�*�`�N����� @_����ҟ|���&� �6�8�J���n����� ȯگ�����"��F��0�  l�p� �p���p��$TB�JOP_GRP �2(8���  ?�p�	�����*���@���@�� 0��  �� � � � ��p� @�l���	 �BL �  �Cр D�����<��E�A�S�<��B$�����@��?�33C�*���8œϞ�� �2�T�����;�2��t��@��?���zӌ�-�kA�>�Ⱥ�� �����l�>�~�a�s��;��pA�?��ff@&ff?�#ff�ϵ�8� ��L����}������:v,����?L~�}ѡ�D�H��5�;�M�@�33`�����>��|օ���8���`ự�	�D"��������`��r�|���"�9������g�v��x��� �������������� 0(V�b������p�C��p�	���	V3�.0�	lr2d��*b��k�p�{ E8� �EJ� E\� �En@ E��E��� E�� E��� E�� E��h E�H E��0 E� EϾ��� E���� E�x E��X F��D��  D�` E��P E�$��0�;�G�R��^p Ek�ui������(��� E�����?X 9�IR4! �H%�
z�`/r"�p�v#Ѭ߱/��E?STPARSI d�쵰��HR� ABL�E 1+��J p��(�' �k)�'��(�(o�w��'	��(
�(�(5p���(�(�(K!�#RDI�/��??(?:?L?^5�4O�?�;�? �?O O2N�"S�?�� �:�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo���@ �O��7�isO�O�O�O U?g?y?�?�?�8�"pb�NUM  8�U����x� J �K �"_CFG �,Y{s�@��IM?EBF_TT�!u8��� �vVERI#�az�v�sR 1-�+O 8mp�k�2� ;��o  �� �,�>�P�b�t����� ����Ώ�����(� :���^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�{�V�h� ��������¿Կ���H
��"�q_Sq�v@�u�� MI_CHA�N�w �u u�DB'GLV���u�u�!�x�ETHERADW ?�%���v ��������(x�R�OUT�p!WJ!�*�H��SNMA�SK���s��255.��N�ߖߨ�N�� OOLOFS_�DI� BŪ�OR�QCTRL .�{>Cw/&�T�J�\� n����������� ���"�4�F�X�j�z���������#PE_�DETAI����P�GL_CONFI�G 4Yyiq���/cell/$�CID$/grp1��;M_q�9C�߮���� �,>Pbt� �����/�� :/L/^/p/�/�/#/�/ �/�/�/ ??�/6?H? Z?l?~?�??1?�?�? �?�?O O�n}�?VO hOzO�O�O�Oq���O�M��?__1_C_U_ g_�?�_�_�_�_�_�_ t_	oo-o?oQocouo o�o�o�o�o�o�o�o );M_q � �������%� 7�I�[�m������� Ǐُ�����!�3�E� W�i�{������ß՟ ������/�A�S�e� w��������ѯ������ �Us�er View �)	}}1234567890J�\�n����������5�	̿��0�2=���� �2�@D�V�h�ǿٿ7�3� �����������o�1�߾4��j�|ߎߠ߲���#���߾5Y��0�B�T�f�x��ߙ�߾6 ���������,���M�߾7��������� ����?�߾8u�: L^p������� lCamera;�1� 0BT2BE�~ ��H�����//�  ���f/ x/�/�/�/�/g�/�/ ?S/,?>?P?b?t?�?�����?�?�?�? OO,O�/PObOtO�? �O�O�O�O�O�O�?�7 XىO>_P_b_t_�_�_ ?O�_�_�_+_oo(o :oLo^o_�72+�_�o �o�o�o�o�_*< N�or����� so���a�(�:�L� ^�p��������܏ � ��$�6���7t� ͏��������ʟܟ��  ��$�o�H�Z�l�~� ����I��7(	9�� � �$�6�H��l�~��� ۯ��ƿؿ���ϵ�ǧ9��O�a�sυϗ� ��P������Ϙ��'�@9�K�]�o߁�
	�0߼��������� ��:�L�^�߂��� ������ߕ�� ��� 5�G�Y�k�}���6�� ����"���1C U���I+����� �����1C� gy����h�� �;X//1/C/U/g/ �/�/�/��/�/�/ 	??-?��![�/y? �?�?�?�?�?z/�?	O Of??OQOcOuO�O�O @?��k0O�O�O	__ -_?_�?c_u_�_�O�_ �_�_�_�_o�O��{ �_Qocouo�o�o�oR_ �o�o�o>o);Mx_qm  i ���������0�B�T�f�    v~������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ�ؿj�  
`( � �p( 	 ���B�0�f�T� ��xϚϜϮ���������,���� � �oq߃ߕ������� ����c`�=�O�a� �߅��������&� ��'�n�K�]�o��� ������������4� #5GYk����� ����1 C�gy���� ���	/P-/?/Q/ �u/�/�/�/�/�// (/??)?p/M?_?q? �?�?�?�/�?�?�?6? O%O7OIO[OmO�?�O �O�O�?�O�O�O_!_ 3_zO�Oi_{_�_�O�_ �_�_�_�_oR_/oAo So�_wo�o�o�o�o�o o�o`o=Oa s���o�o��� 8�'�9�K�]�o�� �������ۏ���� #�5�|�Y�k�}�ď�����şן���B�"�@� �*�<�N���$����+frh�:\tpgl\r�obots\lr�m200id��_�mate_��.xml
���Ưد����� �2�D�V�F��� `���������Ϳ߿� ��'�9�K�b�\ρ� �ϥϷ���������� #�5�G�^�X�}ߏߡ� ������������1� C�Z�T�y������ ������	��-�?�V� P�u������������� ��);R�Lq ������� %7NHm� ������/!/�3/E.g��� |$�r�<< p� ?�E+�/E/�/�/ �/�/�/?�/?<?"? 4?V?�?j?�?�?�?�?��?�?�?
O8OF���$TPGL_OUTPUT 7P��P� h  tE�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo�'otEh �=@2345678901Lo ^opo�o�o�o�cF�Io �o�o�o/�o3@ew���Ez}� ����'���]� o���������O�ŏ� ���#�5�͏C�k�}� ������K�]����� �1�C�۟Q�y����� ����Y�ϯ��	��-� ?�ׯ�u��������� Ͽg�ݿ��)�;�M� �[σϕϧϹ���c� u���%�7�I�[��� iߑߣߵ�����q��߀�!�3�E�W���HA} c!�������������@j/�.�p* ( 	 1oc�Q��� u��������������� )M;q_�� �����7 %GI[��?f�f &��-�#/ 5//Y/k/9j��/�/ H/�/�/�/�/?,?�/ 0?b?�/N?�?�?�?�? �?>?�?O�?OLO^O 8O�O�O�?|O�O�OvO  __�O_H_�O�O~_ �_*_�_�_�_�_�_o l_2oDo�_0ozoTofo �o�o o�o�o�o�o. @dv�o^�� X����*��� `�r����������ޏ <�N��&���2�\�6� H��������ڟt�Ɵ �"���F�X���@��� (�z�į֯�����j� ��B�T��x���d��� ���0���Ϣ��>� �*�tφ�俪ϼ�Vπ��������(�:��)�WGL1.XM�L��o��$TPOFF_LIM �|���}��N_SV��  �����P_MON7 8������2y�STRT?CHK 9�������VTCOM�PAT��6��VW�VAR :��\Y�� � q�������_DE�FPROG %���%MAIN� DT-��u�_D?ISPLAY�������INST_MSwK  �� ��?INUSER,����LCK5���QUI�CKMENY���S7CREx��7�?tpsc��5�Г���ҩ�_��ST�*��RACE_C_FG ;��Y�u��	z�
?���?HNL 2<��`� ��L^p�������
��IT�EM 2=8 ��%$12345�678901 � =<)Oai G !ow��3 �z��A//w )/��v/��/��/ �/M/=/O/a/{/�/�/ �/U?{?�?�/�??'? 9?�?]?	O/OAO�?MO �?�?�?qO�O#O�O�O YO_}O�OX_�Os_�O �_�__�_1_�_og_ 'o�_7o]ooo�_{o�_ 	oo�o?o�o#�o G�o�o�oSk� �;�_q:��U� �y�������%�� I�	�m��?�ŏ��Ǐ ُ���w�!�͟�� i�)�������+�՟�� �����ůA�S�e�� 7���[�m�ѯy���� п+��O��!υ�7� ������߿��ϯ��� ��K���oρϓ�߷� c߉ߛ��Ͽ�#�5�G� ����}�=�O��[��� �߲����1����g�����f���S��>|k��  ��k� ����
 ���������UoD1:\&��}��R_GRP 1?�� 	 @��q�m��������  ��&J5nY?�  ������� /�//'/]/K/�/�o/�/�/�/�/�/�/	�9�?%?{�SCBw 2@�� t q?�?�?�?�?�?�?�?�Oq�UTORIAL A��LOv��V_CONFIG B����	�O�[MOUTPUT �C���@�� �O�O__1_C_U_g_ y_�_�_�_�_�_�A�O �_oo1oCoUogoyo �o�o�o�o�o�_�o	 -?Qcu�� ����o���)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ���������'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���������� �O�E�O'�9�K�]�o� ���������������� ��#5GYk}� ������ 1CUgy��� ����	/-/?/ Q/c/u/�/�/�/�/�/ �/�/?/)?;?M?_? q?�?�?�?�?�?�?�? O?%O7OIO[OmOO �O�O�O�O�O�O�O_  O3_E_W_i_{_�_�_ �_�_�_�_�_o_/o AoSoeowo�o�o�o�o �o�o�oo+=O as������ ���&9�K�]�o� ��������ɏۏ���|������0� B�,��m�������� ǟٟ����!�3�E� W�i��������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sτ� �ϩϻ��������� '�9�K�]�o߀ϓߥ� �����������#�5� G�Y�k�}�ߡ���� ��������1�C�U� g�y������������ ��	-?Qcu �������� );M_q�� �����//%/ 7/I/[/m//��/�/ �/�/�/�/?!?3?E?�W?i?{?�;�$TX�_SCREEN �1DD��,��}ipnl�/�0gen.htm�?�?�?OO%O���Panel �setup)L}��)OjO|O�O�O�O�O XONO�O__1_C_U_ �Oy_�O�_�_�_�_�_ �_n_�_-o?oQocouo �o�_,o"o�o�o�o )�oM�oq�� ���BT��%� 7�I�[�� ������ Ǐُ���t�!���E��W�i�{�������>U�ALRM_MSG� ?�9��0  ���*��5�(�Y�L� }�p�������ׯʯ�����ӕSEV  ��Q�ђEC�FG F�5�1  �%@� � A��   B��$
  ��#�5�� ƿؿ���� �2�D��V�h�v�]�GRP �2Gg� 0�&	� ����ӐI_B�BL_NOTE �Hg�T�G�l�"�0�!s�~��DEFPROݐ=%� (%�:� � (�a�L߅�pߩߔ� �߸������'��K����FKEYDAT�A 1I�9��p v��&�ϰ���0��������,(�+���$(POINT�  ]3�5���NC�EL_����NDI�RECT���� EXT STEP���6�TOUCHU����ORE INFOOaH �l�������9 ]o ���/frh/�gui/whit�ehome.pn�gp������}�point��*/</N/`/r/&  �FRH/FCGT�P/wzcancel/�/�/�/�/�/��#�indirec/4?F?X?j?|?�/� nex#?�?�?�?��? O$�touchup�?<ONO`O�rO�O$�arwrg�?�O�O�O�O_ �8#_5_G_Y_k_}_�_ _�_�_�_�_�_o�_ 1oCoUogoyo�oo�o �o�o�o�o	�o? Qcu��(�� �����;�M�_� q�������~��ӏ� ��	��-�4�Q�c�u� ������:�ϟ��� �)���;�_�q����� ����H�ݯ���%� 7�Ư[�m�������� D�ǿ����!�3�E� Կi�{ύϟϱ���R� ������/�A���S� w߉ߛ߭߿���`��� ��+�=�O���s�� ������\����� '�9�K�]��������з�����v���>����# 5WiC,U� M������ <N5rY��� ���/�&//J/ 1/n/�/g/�/�/�/�/ ���/?"?4?F?X?g� |?�?�?�?�?�?�?w? OO0OBOTOfO�?�O �O�O�O�O�OsO__ ,_>_P_b_t__�_�_ �_�_�_�_�_o(o:o Lo^opo�_�o�o�o�o �o�o �o$6HZ l~����� �� �2�D�V�h�z� �����ԏ���
� ��.�@�R�d�v���� ����П������/ <�N�`�r��������� ̯ޯ���&���J� \�n�������3�ȿڿ ����"ϱ�F�X�j� |ώϠϲ�A������� ��0߿�T�f�xߊ� �߮�=��������� ,�>���b�t���� ��K�������(�:� ��^�p����������� Y��� $6H�� l~����U��� 2DV-��X�-�������}���,�/
/�/.//R/d/ K/�/o/�/�/�/�/�/ ??�/<?#?`?r?Y? �?}?�?�?�?�?�?O �?8OJO)�nO�O�O�O �O�O��O�O_"_4_ F_X_�O|_�_�_�_�_ �_e_�_oo0oBoTo �_xo�o�o�o�o�o�o so,>Pb�o ������o� �(�:�L�^�p���� ����ʏ܏�}��$� 6�H�Z�l��������� Ɵ؟����� �2�D� V�h�z�	�����¯ԯ ������.�@�R�d� v���_O����п��� ��*�<�N�`�rτ� ��%Ϻ��������� ��8�J�\�n߀ߒ�!� �����������"�� F�X�j�|���/��� ����������B�T� f�x�������=����� ��,��Pbt ���9��� (:�^p�� ��G�� //$/ 6/�Z/l/~/�/�/�/��/���+�������/?=�/7?I?#6,5Oz?-O�? �?�?�?�?�?�?O.O ORO9OvO�OoO�O�O �O�O�O_�O*__N_ `_G_�_k_�_�_���_ �_oo&o8oG/\ono �o�o�o�o�oWo�o�o "4F�oj|� ���S���� 0�B�T��x������� ��ҏa�����,�>� P�ߏt���������Ο ��o���(�:�L�^� ퟂ�������ʯܯk�  ��$�6�H�Z�l��� ������ƿؿ�y��  �2�D�V�h����Ϟ� �����������_�.� @�R�d�v�}Ϛ߬߾� ��������*�<�N� `�r��������� �����&�8�J�\�n� ����!����������� ��4FXj|� ����� �BTfx��+ ����//�>/ P/b/t/�/�/�/9/�/ �/�/??(?�/L?^? p?�?�?�?5?�?�?�?� OO$O6O�8K}�����aO@sO�M]O�O�O�F,�_ �O�__�O2_D_+_h_ O_�_�_�_�_�_�_�_ �_oo@oRo9ovo]o �o�o�o�o�o�o�o *	�N`r��� �?�����&�8� �\�n���������E� ڏ����"�4�ÏX� j�|�������ğS�� ����0�B�џf�x� ��������O����� �,�>�P�߯t����� ����ο]����(� :�L�ۿpςϔϦϸ� ����k� ��$�6�H� Z���~ߐߢߴ����� g���� �2�D�V�h� ?������������ 
��.�@�R�d�v�� �������������� *<N`r�� �����&8 J\n���� ����"/4/F/X/ j/|/�//�/�/�/�/ �/?�/0?B?T?f?x? �??�?�?�?�?�?O O�?>OPObOtO�O�O 'O�O�O�O�O__�O :_L_^_p_�_�_�_}���[�}�����_�_�]�_o)of,Zo~oeo�o �o�o�o�o�o�o2 VhO�s�� ���
��.�@�'� d�K�����yﾏЏ� ���'_<�N�`�r� ������7�̟ޟ�� �&���J�\�n����� ��3�ȯگ����"� 4�ïX�j�|������� A�ֿ�����0Ͽ� T�f�xϊϜϮ���O� ������,�>���b� t߆ߘߪ߼�K����� ��(�:�L���p�� ������Y��� �� $�6�H���l�~����� ���������� 2 DV]�z���� ��u
.@R d������� q//*/</N/`/r/ /�/�/�/�/�/�// ?&?8?J?\?n?�/�? �?�?�?�?�?�?�?"O 4OFOXOjO|OO�O�O �O�O�O�O�O_0_B_ T_f_x_�__�_�_�_ �_�_o�_,o>oPobo to�oo�o�o�o�o�oh��{������ASe}=��sv,���}� ���$��H�/�l� ~�e�����Ə؏���� � �2��V�=�z�a� ������ԟ����
��� .�@�R�d�v����o�� ��Я�������<� N�`�r�����%���̿ ޿��ϣ�8�J�\� nπϒϤ�3������� ���"߱�F�X�j�|� �ߠ�/���������� �0��T�f�x��� ��=���������,� ��P�b�t��������� K�����(:�� ^p����G� � $6H�l ~������� / /2/D/V/�z/�/ �/�/�/�/c/�/
?? .?@?R?�/v?�?�?�? �?�?�?q?OO*O<O NO`O�?�O�O�O�O�O �OmO__&_8_J_\_ n_�O�_�_�_�_�_�_ {_o"o4oFoXojo�_ �o�o�o�o�o�o�o�o 0BTfx� �������,�@>�P�b�t���]����]������ÏՍ����	��, ��:��^�E�����{� ����ܟ�՟���6� H�/�l�S�������Ư ���ѯ� ��D�+� h�z�Y����¿Կ� ����.�@�R�d�v� ��ϬϾ�������� ��*�<�N�`�r߄�� �ߺ���������� 8�J�\�n���!�� �����������4�F� X�j�|�����/����� ������BTf x��+���� ,�Pbt� ��9���// (/�L/^/p/�/�/�/ �/���/�/ ??$?6? =/Z?l?~?�?�?�?�? U?�?�?O O2ODO�? hOzO�O�O�O�OQO�O �O
__._@_R_�Ov_ �_�_�_�_�___�_o o*o<oNo�_ro�o�o �o�o�o�omo& 8J\�o���� ��i��"�4�F� X�j��������ď֏ �w���0�B�T�f� ����������ҟ����� ���� ���!�3�E��g�y�S�,e���]�ί�� ���(��L�^�E� ��i�������ܿÿ � ���6��Z�A�~ϐ� wϴϛ������/� � 2�D�V�h�w��ߞ߰� �������߇��.�@� R�d�v������� ������*�<�N�`� r�������������� ��&8J\n� ������ �4FXj|� �����/�0/ B/T/f/x/�/�/+/�/ �/�/�/??�/>?P? b?t?�?�?'?�?�?�? �?OO(O��LO^OpO �O�O�O�?�O�O�O _ _$_6_�OZ_l_~_�_ �_�_C_�_�_�_o o 2o�_Vohozo�o�o�o �oQo�o�o
.@ �odv����M ����*�<�N�� r���������̏[��� ��&�8�J�ُn��� ������ȟڟi���� "�4�F�X��|����� ��į֯e�����0��B�T�f��$UI_�INUSER  �������  g��k�_MENHIS�T 1J���  (���?@(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1���+�=�Oπ9)��631Ϝ�������a�s�edi=t��MAIN�� �82�D�V� �'��v΁2ϡ߳������� ����%�7�I�[��� ��������h��� �!�3�E�W���h���@������������{� ۱{�*<N`r u������� &8J\n� �������"/ 4/F/X/j/|//�/�/ �/�/�/�/�/�/0?B? T?f?x?�??�?�?�? �?�?O��>OPObO tO�O�O�?�O�O�O�O __�O:_L_^_p_�_ �_�_5_�_�_�_ oo $o�_HoZolo~o�o�o 1o�o�o�o�o 2 �oVhz���? ���
��.�O+O d�v����������� ���*�<�ˏ`�r� ��������̟[��� �&�8�J�ٟn����� ����ȯW�����"� 4�F�X��|������� Ŀֿe�����0�B� T�?�Q��ϜϮ����� �����,�>�P�b� ��ߘߪ߼������� ���(�:�L�^�p��� ����������}�� $�6�H�Z�l�~���� ������������ 2�DVhze���$�UI_PANED�ATA 1L����� � 	�}/f�rh/gui�d�ev0.stm �M?connid�=0 height=100&_� �ice=TP&_�lines=15�&_column�s=4� font�=24&_page=whole� ��h�)prim/X  }[�0���� )�� �#/
/G/Y/@/}/d/ �/�/�/�/�/�/?�/�1?h��� �    ��in?�?�?�?�? �??�?_O"O4OFO XOjO�?�O�O�O�O�O �O�O�O__B_T_;_�x___�_�_�_�_E7  � �U�Oo$o6oHo Zolo�_�oO�o�o�o �o�ouo2D+h O������� 
���@�'�d�v��_ �_����Џ���Y� *��oN�`�r������� ��!�ޟş��&�8� �\�C�����y����� گ�ӯ�����F�X� j�|������ĿֿI� ����0�B�Tϻ�x� _ϜϮϕ��Ϲ���� ��,��P�b�I߆�m� ���/������(� :�L��p�㿔��� ������U��$��H� /�l�~�e��������� ������ DV�� �ߌ�����9 
}�.@Rdv� �����// �</#/`/r/Y/�/}/ �/�/�/�/cu&?8? J?\?n?�?�/�?�?) �?�?�?O"O4O�?XO ?O|O�OuO�O�O�O�O �O_�O0_B_)_f_M_�_�/?}��_�_�_�_
oo.o)�_So�5 Boo�o�o�o�o�o@o �o�o!W>{ b���������/��83;�$U�I_POSTYP�E  5?� 	 ;����a�QUICKME/N  p�����c�RESTORE� 1M5�  �*default�;�SINGLE~ԍPRIMԏ�mmenupage,23,1<� n�������G���П� ������<�N�`�r� ���"������ϯ�� 
��.�@��d�v��� ����O�п����� ï%�7�Iϻ��ϖϨ� ����o�����&�8� J���n߀ߒߤ߶�a� ������Y�"�4�F�X� j���������y� ����0�B�����a� s������������ ��,>Pbt�������SCR�E��?���u1sc�u2�!3!4!5!6�!7!8!�TATl�� ă5Y��USERTL#ks+�4�U5�6�7�8��a�NDO_CFG� Np��P�Qa�O�P_CRM5  ��U&a�PDd���Non�e���_INFOW 1O5f 0%��/�8o/�/�/ �/�/�/
??�/@?#? d?v?Y?�?�?�?�?���S!OFFSET Rp�j!�?��� �!O3OEOWO�O{O�O �O�O�OO�O___ J_A_S_�_w_�_�_�Kŏ�]�_
o
�_/o�8UFRAM%�/P!�RTOL_ABRqTSoN#kbENBto~ehGRP 1S�����Cz  A� �c�a��o�o�o�oB"v,>cj��U�h�#!�kMSK  h�ef!�kNPa%^)��%�_��e_EV�Ns`�t&�v�2�T�;
 h#!�UEVs`!td�:\event_�user\�7�C�7<�o� Fq�/�S�P5�:�spot�weldl�!CA6��r���#�t!� K�	�>��q��-�� q���Q�c�ܟ�� ��� ��ϟH��l��)�_� ����د����˯ �� D���z�%�����[��m�濑�
ϵ�Ǻ�W�RK 2U�a8�nπ� \ϥϷ� ���������#���G� Y�4�}ߏ�j߳��ߠ� �������1��B�g��y��$VARS__CONFI�V�;� FP����C�MR�b2\�;�xy� 	$ ��0�1: SC130EF2 *�	�����X�ȸp�  �#!?�p@pp:"p�z� o]�g���������������`�uA�����,� B���G�K��l�� �_������ �2�hSe��Q����IA_W�OF�]^-˶,�		�Q;%/+'G��P �> ���RT�WINURL ?5�������/��/�/�/�/�/�SI�ONTMOU� ���%�^Sۿ��S۵@�a� FR:\�#\�DATA؏  �� UD166wLOGC?  \9�EXh?'q' ?B@ ���2{1�U��?{1�?�?θ �� n6  �������2zt�`�F��  =����BA��?@|=TRACIN�?AQB�d�CpBEFF/B�0�(��_� (��I�M ��O�O�O__P_>_ t_b_|_�_�_�_�_�_.�(_GE3`�/C��
�`'p4b
g�0R�E!0a�i���LE�Xdb����1-e��/VMPHASE'  ���C ���RTD_FILT�ER 2c� �&��T��o+ =Oas�����o ������1�C��U�g��)SHIFTMENU 1d�K/
 <�<%�?ŏ2����ɏ�ُ� 8��!�n�E�W�}���������ß՟"����	LIVE/SN�A��%vsflsiv�n4���#� SETU��W�menum�r��ѯ��"��3e`+|�MO�3ftn�z��ZD��gQm˳<�A�P��$WAITDINEND8L!�k�OK  �醼 :r��S����TIM5���Gr�͔��%˴��ӿ�򿆸RELE�a5��k��/<6m�_ACTJ�4�t !��_?1 h���%�5߅���RD�IS����$X�VRnaitn�$oZABC��1jQk' ,�@�2=��-�ZIP2kQo����)���MPC?F_G 1l��l!a0L"��q�7�MP��am����P�������`�*�  4�Y��G�4/���G�Y�Ǵ��K�y5�����H�D�b���_�B��B�0�Q��5�(>����<�ȴ0+&���=I?�j�\����&?���|���&?���{� ?�.��8�}���p9��������C²��B���j�r�7�5B��³ a´ 'Gl�PJ\r� �������6��.�ȇ�J�p`n��_C_YLIND�aoR�� �p6 ,(  *o�w3l���� ��// '.iJ/�n/U/g/�/ ��/�/�///?�/�/ F?-?j?Q?�/�?�?r�Cp*� �g� �?L^���6O!OZO?Ih�?�O?G��AA�=�SPHERE 2qO�?�OT?�O_ �O:_�?�Op_�_�/�_ E_+_�_�_ o�_Y_6o Ho�_�_~o�_�o�o�o��oo�o ��ZZ�� ��