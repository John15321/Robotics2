��   t�A��*SYST�EM*��V9.1�035 7/1�9/2017 �A   ����DMR_GRP�_T  � �$MA��R_D�ONE  $�OT_MINUS�   	GPyLN8COUNP �T REF>wP�OOtlTpB�CKLSH_SI�GoSEACHMsST>pSPC�
��MOVB RAD�APT_INERzP �FRIC�
_COL_P M�
�GRAV��� HsIS��DSP?��HIFT_ER[RO�  �NA�pMCHY SwARM_PARA#w d7ANGC �M2pCLDE|�CALIB� �DB$GEARz�2� RING���<$1_8k����CLC.o � �AXO � $PS_�T�I���TIME� mJ� _CM�D�T"FB�VE}Lg'CL_OVj�~ FRMZ�$DE��DX�$NAM {%�CURL� �kWu�mTCK��%�FMS*��REM_LIF��u�(�*'$��)_0�*_�����#(6+~ K"lPCgCOMi�FBk yMV0�MAL_�#EC�S�P!3"7DTY?R_@"�5��#�1END�4���C1  P�L~ + ��S�TA�#TRQ_MH��� K"FS� �)HY'J� GI4JI�BJIPD��$�A�SS  �����A�����@V�ERSI� �G  �ӞA?IRTUAL�O�A�' 1 �H � �� 	 ��_�O4__X_?_ |_g_y_�_�Z�@�_�\ИA�_�\�@� O������A�Y`���+�_Do�_	l�boto�o�o�o�o8k �o�b�o-Q���dAz����=L3�ͩ�?����@���(�:�L�^� p���������ʏ܏/ �E����5��D  2if�x����������ҟ������< U�2�D�V�h�z��������¯ԯ������@���$�$ 1�L��?qN�f�N��O�M���Eڻ� D�F@2~@�0��@+��?���s)���:b�7^j63}B�p����������еA�: ϯ: Ƚ8�J�п]�Hρ�l���Ϸ��LL�Kp�������� ��� ��ߘ�9�$�]�o����%R�345678901�ߗԼ���%� ��!������.�K��� N�`���6��ߐ��� ������@��#�v��� V�D�z�h�������� *�<�����
@.d ��������N� �*�Qc� ������F/ j|��J/�/n/�/ �/�/0/B/?�/4? "?D?j?�/�?�?�/X? �?�?�?�?O0O�?WO �?�?6OO�O�O�O�O :OLO_pO�OP_�Ot_ b_�_�_ _�_�_6_�_ oo:o(o^opo�_�o �_�_voHo�o �o$ zo�o]�o�o�� ���@�#�v� V�D�z�h������׏ *�<�����
�@�.�d� ��̏�����ПN��� ��*���Q�c���� ��������ޯ�F�� j�|���ȯJ���n���රű�ݿ0��$P�LCL_GRP �1 ��� DT�?�  &�8�X�[�T��j� �ώ��ϲ�������!� �E�W�