��   �A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����BIN_C�FG_T   �X 	$ENTR�IES  $�Q0FP?NG1�F1O2F2OP�z ?CNETG����DHCP_C�TRL.  0{ 7 ABLE? �$IPUS�R�ETRAT�$SETHOST��NSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!� FT� =@� LOG_8	,�CMO>$DN�LD_FILTE�R�SUBDIR'CAPC����8 .. 4� H{ADDRTYP�=H NGTH��f��z +LSq� D $RO�BOTIG �PE�ER�� MASKn�MRU~OMG�DEV��PIN�FO�  �$$$TI ���RCM+?T A$( /�QSIZ�!S~� TATUS_%�$MAILSER�V $PLAN~� <$LIN�<$CLU��<�$TO�P$CC�&FR�&YJEC�|!Z%ENB ^� ALAR:!B��TP,�#,V8 S���$VAR�)M��ON�&���&APPL�&PA� �%�N�'POR�Y#_�!>�"ALERT�&i2URL }Z3�ATTAC��0ERR_THROU3�US�9H!�8� CH�- c%�4MAX?W�S_|1��1MOD��1I�  �1�o (�1PWD � � LA��0�N�D�1TRYFDE�LA-C�0G'AERcSI��1Q'ROBICLK_HM 0Q'� �XML+ 3SGF�RMU3T� !OU�U3 G_�-COP 1�F33�AQ'C[2�%�B_AU�� 9 R��!UPDb&PC�OU{!�CFO ?2 
$V*W��@c%ACC_HYQS�NA�UMMY1�oW2?��RDM�* $DISL��SN,#	3 ��	o!�"%"_W�I�CTZ_IND9E�3�POFF� ~UR�YD��S�  
 t Z!KRT�0N�(cD�.)bHOUU#E%A/f�Va>fVaMfLOCAܗ #$NS0H_[HE���@I��/  d�PARP�H&�_IPF�W�_* O�F�PQF�AsD90�VHO_�� 5R42PS�a?�wTEL� P����90WORjAXQE� LV�O#�FS1�ICEد[p� �$�c  ����zq��
���
op�PS�Axw�# �i�qIz0ALw�q'0 �x+
���F�����p��r�u�$� 2�{���r#���� �}��!�qi�����$� _FLTRs  �y�p ��������}�$��}2}��bSHARV� 1�y Pe���t
�G�6�k�.� ��R���v������� П1���U��y�<��� `�r�ӯ�������ޯ ?���u�8���\��� ��ῤ�ڿ��;��� _�"σ�FϏ�jϸ��� �����%���I��m� 0�Bߣ�f��ߊ��߮� �����E��i�,�� P��t����������/���z _LUA1���x!1.j�0�8���i�1z���2�55.��q�����uh�2o��������������3����^ 1C��4_���  ������5���@N�!3��6O����u�������QJ���� ��(�� Q� '��<a/�/�/{/�/@�/�/�/?&?��P? V?h?z?9?�?�?�?�? �?�?
OO��?����ufOQL
ZDT Status�?�uO�O�O�O��}i�RConnect�: irc�D//alert�N&_8_ J_\_�G�O�_�_�_�_(�_�_���sP 2ـd���_o1oCoUo goyo�o�o�o�o�o�o��o�s$$c962�b37a-1ac�0-eb2a-f�1c7-8c6e�b5f01a8c  (y_J�On�H�����ـP(�X"�rZJ�u3 �v[C] )�,$e"�ـ[� �M�4�q�X�~����� ˏ�����%��I��0�B��f���������w�W�8 DM_�=!W�G�SNT-P�	�%��-�����������K�4#��USTOM' 
�F��W � �3$TCPIP��XHO%S"���ELO�W�T!�E�H!Tb����rj3_tp�dQO \��!KCL�������v!CRTY�G����O"(�!CON�S�� ��ib_Osmon����