��  	w^�A��*SYST�EM*��V9.1�0185 12�/11/2019� A  �����AAVM_�WRK_T  �� $EXP�OSURE  �$CAMCLB�DAT@ $PS_TRGVT��$X aH]ZgDISfWg�PgRgLENS_CENT_X��YgyORf  � $CMP_G�C_�UTNUM�APRE_MASwT_C� 	��GRV_M{$�NEW��	ST�AT_RUNAR�ES_ER�VTSCP6� aTCb32:dXSM�p&&�#END!�ORGBK!SMp��3!UPD�O�ABS; � P/ �  $P�ARA�  ����AIO_wCNV� l� �RAC�LO�M�OD_TYP@F+IR�HAL�>#�IN_OU�FA�C� gINTER�CEPfBI�I�Z@!LRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CESI0�!H1�!"PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W� @V�R!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2 � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1 UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t�cbMO� �sE 	� [M�s��2�wREV�BILF��!XI� %�R 7 � OD}`j��$NO`M��i`�x�/�"u�� ����^���@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQC���a_EDu �O � C2��`�S�p�4%$l �t'$OP�@QB�qy��_OK���0, P_�C� y��dh�U �`LACI�!�a���<� FqCOMM� �0$D��ϑ�@�pX���ORgf�BIG�ALLOW� �(KD2�2�@VAaR5�d!�A}#BL[@S � ,KJqM�rH`S�pZ@M_O]�z���CFd X�0GR@��=M�NFLI���;@UIRE�84�"�� SWIT=$/0_uNo`S�"CF_��G� �0WA�RNMxp�d�%`L�I�V`NST� C�OR-rFLT�R�TRAT T|�`� $ACCq�S�� X�r$OR�I�.&ӧRT�`_�SFg��HGV0I��p�T��PA�I
��T��0��� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8� �
���x@�2� @� TRQB��$%f��ր����c_U���� COc <� ����Ȩx3�2��LLECM�}-�MULTIV4��"$��A
2FS�I�LDD��c� DET}_1b  4� STY2�b4�=@��)24��e`DԼ� |9$��.p��6�aI`�* \�TO�:�E��EXT����p���B�ў22f�,E��@��1b�.'�B ��G�Q� �"Q�/%�a��X� %�?sdaD�U� Sҟ؈;A�Ɨ�M�� �� CՋO�! L@�0a�� X׻pAβ�$JOBB���� � ��IGO�" d Ӏ�����X�-'x���0G�ҧ����_M��b�# tӀF� �CNG�AiBA� ϑ�� !���/1��À�0����R0P/p����$
�|��BqF]��
2J]�_RN��C�`J`�e�J?�D/5C�	�ӧ��@���P�O3л!% \��0RO�6� �IyT�s� NOM_8p�n#�c ���T5U�@P� � ��E&+P��� ӨP�	ݭ��RAx@n �3�<A���
$TF3%#KD3
T��wpU�1�3�}�%mHrzT1�E���ޣ�#�ݤ�%ߢQlYNT|�"� DBGDE�!3'D�]�PU���@0t����"��AX��"�uTAI2sBUF8ۆ;%�1( ��P&�V`PI84'mP��'M�(M�)B �&F>�'SIMQS�@ZwKEE3PAT��zЙ8"�"԰��Cb��)S�0��`JB���ľaDECg:� g5�e�����* �U�CHNS_EMPͲG$G��7�_�<�c;�1_FP)�TC�6S���5�`%��4�} ��V����W��JR����SEGFRAq�O�� #P�T_LIN�KCP�VF����C$+ ���ckBZ��PBzr��|�@6,` +� Ԧ��A�0��Ad0o`�Ar�D���Id1SIZh���	T�FT�C�Z1Y�ARSm��CP@�'�Ic\1@cX�0<@Lp����0�VCRCߥ�sCC���U1@�X�1��2�Mpq�U�1`��X�Q�UDݤأiC k�p��
DK`݀f��RhEVRf �Fha_
	EF�0N�f�Pd1��&h��5�jC}�+��VSCA[��A��f�B�4��-�	<�ׇMARG���"a�F@@���1DcQ�rN�0LEW�-��R��P<��o�l��RɄ.� ����ǯ��� 5ڡR�`HANC��$LG5��a��Ӑ��ـF��Ae����0RYr�3
����
��@ �RA��
�AZ��0Q�N`�O��FCT��sp�F��R�0\P0b ADI��O�� +���+���&���5�5Є���S[�g���BMPUD(PY�1��GAESCPjc��W���N  SuU0ۑU:�/)�TIT'q<��b�%ECA:!�!ERRLd��0�&Q��OR�B$��������?$RUN_O��SYS��4������Nu�REV�c� ��OPXWO�P�10�$SKo�"vЂ��T�pTRL�2 �C AC����%�m�&U DJ�p�_p�!�A�ǀM�PL�A�_2WA��j�E��D�!w�!�BhO�UOMMY9����1Л / DB[��3����!PR�Qe�f�qDٱ9��4 ж�$r�$ Q��Lة5�z�����6�z��PC�7*�<�EN5EC0Tq8I�����RECOR$�9�H m��4$L��5$أ�"E�`��R@��VA��_Dց�� ROS) �"SK �����I�=�א���PA��JVBETU�RN���SMR(�U�) #�CRʰEWMzDB0GNALV ��"$LA� [�*�6$P-�7$P�v�s�8o�!�PC��#�DO^@-�Ŵ����R˶GO_AW��ܱMOz��p��d�DCSS_CN4�YO�:��T��0L���ID�T�2��2�N��O@�J���v`Iְ ; P7 $>�RB�B���PI�POl�I_#BY��vЅ�TVR���HNDG$�< �H�`�1a�@cS��DSBLI��s���0Z}�p��LS$�=�Ҙ0� ��FB�FEձL�9����5��=>D�$DO�1�C�pMC�0q��4��9�RH��W��K4ELE�ur������SLAVr?xBIANS ���#����_R@P�@\`�pS�}��l�}�l�{u��[!e��ے�I���B��9W��D�NTV�#�sVE�$��SKI�lA4;3��2UB�1Jp�f�1C�
DSAF7��5��_SV6�EX�CLU-��XrONL�0YY��s�����HI_VՀ�RPWPLYo�RCsH� ��0_M�Q�VORFY_I�.Mms$IOv0��}���1UB���Oj�3LQS����4!�R�:@�P�$��~�AUTOCNE �����.��GCH�D�s��_���3s�AMF��CPe�T!q��р� Ao����_�0  .��NOCtBxB�p	T��A ��z��SG�` C �? 
$CUR8�U� �!" �� T@B���|��ANNUNC�@#���䱐b����()%!��-*I&���tp@��IC�D @�1F
"a��POTX�aӀ����������֠E-M��NIߢE�·"�G� A��$DAY��LOAD`Ԟ��"���5���EFF�_AXI�Fo��%Q�O0�:�_RwTRQV1G D�a��?0�RK3�0S45 2Fz@]w:1a���A0p/1sAH 	0B!�1A�T�2�ûv�DUX��u��CAeBsAIs"�pNS�16�PID�@PWSs�54�AWpV`�V_�0q0>�P�DIAGysAJ� 1$VX��ET	`�UrT��EJ��b{RRf��!�TVE�� SW|AZ�sP��0�:5q0G}P:1O�HP5�1PP|@�SI	R|�{RB�P�2�3%q ZQC �BB��H�^��E`��5q0I��?0��ދURQDW�EMS�B�?UA�p�EjB�TLIFEp[#iP��uRN|QFB�U%!zSFB�a��%"C���Nr��Y'p�FLA�tf& OVڰ�VHE�>�BSUPPO(���uRI�_�T��Q_�X�d�� gZjW�j� g��%!��6�X�Z*�ϡfAY2xhC"��T��DEN�pBE*%!J�� �F_8p�Ax���p�K `QЏCACH�*r�bSCIZ�V�P`�N��oUFFI`� oP�ў�2��6����M;��tL 81 K�EYIMAG �TM��!�^q:�Yv���>��OCVIE�@�q'M �༠L~���;�?��`��р�dN�G0��ST��! �r���t���t� �t0>�pEMAILo���x�!��5FAUL�"�O�r��/���COU����η�T��)AP�< $9�p�S�0�0IT��BUF@�g;��gE�o�e��P	Be�p�C:���:�|�G�SAV��r�[@�b ��@ˇÐ)&P��p����D��_e���� �#OT겮�3Pm ��0�z3�AX�#f x �Xe�C�_G|S
�>�YN_�A��Q E<�Dk�O����BUM�2�PT� F!��$�DI[E�7�����R��$ G���!&�Ǳ����:�9�S����-�&�C_ᰤ�K�$�����RVq���gDSPnv�PCe�IM��\���<�3@�U9��P�] �IP`���A�`[�TH�`�3�O�0T�\�HSȓ>�BSC���`e�V��
��#���*4NV��G;���`Y�e�F|A}�d>���Z��"�SC%Ba��ME�R)�FBCMP�)�ET�� T6LrFU`DUY���R�mb�CDR�ܠ'�6"�f��NO�n!UG0*����%���%)P���C�
ō�\"2��:�o VH *
�L��)� 9���G ���}�Z{� �!{ư!{�1{�6q{�7x�8x�9x�|PzȪ��1��1��1��1���1��1��1��1J��2��2�ˑ�2��U2��2��2��2��U2��2��3��3�ʩ3�˞�3��3��3���3��3��3��4��1EXT6An!W ��߸���V��uş�����`FDR%DXTE�V� .�uR��
�uRREM^@F����BOVM5�*�A�3�TROV3�DTl��S�MXb�IN3�8�PR�"AINDq�cB!
��ɐ}���Ge��C�\�p�UkADO6\�R�IVW�R�BGEA-R5�IObEK#�cDN��1`X� zp`>dCZ_MCMp`uQ� �F�PUR��Y� ,���? ̼P>?o {A?EoE� w����\����Z )QPM��2@RIᵄr�E�TUP2_ [ � q�TDʠ�1p��T�����r�B;AC��\ T�pr�
�)�%w#@ó�TIFI�A����d��@�/PT�B5�FLU=I�t] �@�x;�UR�A���R�БP
��:C_0I�$�]S_?x�J�sCO��"�VRT��>� x$SHO^14 #�ASS�-��U̠��BG_ �!.�!���!��!��FOR�C#�� jDATAZ)A^�rFUZ1��:]#2��LOGh�`�)A_ |��NAVN=�������S��S$VIS�I��SC=�SE�� ��5V� O�1�&1BF�4@�&$�PO� I�A��FMR2��` ���2���6 �!3J�)�CE#��_����_@IT_�Yִ]@M������D�GCLF�EDGDMY�8LD���5�VH���T�M���sa� �v9 T�FS
��tb P��RB��>}�$EX_RAiHBRA1Y�X��RS@3�K�5�F�G&�	5c Y�� ��SW��O0VDEBUG$�A(��GR� opUz�BK�U��O1M� �0POZ0Y�@���E:�@M�LOOM�9QSM�0E������P_E d �P��K�TERM[Ue~dV�ORI֑r`PfdV��SM_㐄�`PgdV� Q �Xh��YUP�ri� -���2d�rS�P�e� G�Z @ELT�O���A�FIG��bZ �A�`�T�Tf�$UFR�$`��aM`ѵ�0OTZg�A�TA��lcNSTאPAT��`�bOPTHJ�ϰE�p8�ذbART؀"ep)�؁���REL�j�SHFTӢ�a��h_�R��̳�V �P$�Wph�1�����t�SHI�`�4Uz � ҁAYLO�� �1��l� ��a}!�ޠERV��Sq�x ��hgא�b �K�u.��KRC��ASY1M���WJ+g�Ⴃ�E��a�y�ұU��א���e@�v�eP���ppE�2vORאML3��GRJQ
4jX"��B0V�`G`�1� HO�6Dk ��aN� ��OCaQ@$OP�$e�i��#����Հ�RY��aOU��c�PTR�e����a�e$PWR��IM��rR_˃�d� �P̛cUD��cSV���֔l� $Hz�!��ADDR��HMQG�b������ ����!1m H��S ���! ��.�畞��ƫ�SEz1�# HS<ܰ
3n $Z À�_D��P�.�PR�M_�"eHTT�P_��H1o (��OBJ� ��$��LEyc��d��p � �睱AKB_��T@S��S����{KRLK�HITCOU� À�! 퀶�����M��SS��v�JQUE?RY_FLA!a���B_WEBSOC��"�HW��a1q��7�INCPUR�!Ou�ˡ�Č������������IO�LNr 8��R�	� $SL2$INPUT_PQ�$�ܸP�# ���SLA�1 sðٿ���s���rNAIOC�F_A5S8Bt$t ��
[�Nq�!]�/a�0ɳ�@ҳUpHY����lïAG�UOP5Eu `X������ā������P������ �����UQ� M�qqgv l�@;sTAkr��A�TI��.�a��Z0S��`PSR�BUZ0ID~0��z���`y�lQ!�u�z`w�"3�f�G��N��Z0>���IRCA���_ x Ĩ��CY�EA{���! ���%�R�`�q<|�8�DAY_��}�NTVA���i��8�eu�i�SCAepi�#CL�������� �qy���ԧb����N_ՀCQ�Ђ�W�rz�O ���������y�G�]�O! 2yG d �q{8P���P�LABzan�\Z0t�UNISb��PITY��"ѳ���IR$6D|R�_URL� �$AL10EN�@�� �P�H�T�T_U� s�Jt�q} X��t�R��" �0�A�D�,J�8F�Lt@�80
K�3
��UJR	5~ ����F|@1w�FgwD^��$J72�O!�/$J8�	7�@\�$��7s�� 8�	�oAPHI@Q�z�Df@J7J8��
L_KE�� o �K��LM���  <��XR�K��� �WATCH�_VA�!pp��F/IELD��y+�&&��� �0paVyp���CT��E��B`��LG���� �!��LG_SIZ����@�3@�O��FD�I��,Q�� ]P����J&3@J& O�J&�J&]PJ&�q�E`1_CM^c�!{@�*h1F��'�$��9(�#r��&@3@�&O��&��'I�(��(,P�&]P�&�RS�I�`  (�PL)N��B�����@ {A�g1��K�u1���L~3t2DAU�5E�AS������2�0GH�����[�BOOܑ��� Cr�[�IaT8��4<`n�RE(Ў�8SCR� ڣs�D�Im�SG`G@RGIPR$D/L�f�քYB$��[�S��Z�W7D[�܉4f�JGM�GMN3CHH�[�FN�F1K�G��IUF�H2pn�HFWD�HHL�ISTP�JV�H�P�H,�0�HRS3YHJ��Kc�C4tS�f�x�kG�YUJ��DjG 3yE�d{��BG�I�`PO�W`Z&ES�"�DOC��v�FEXb�TUI�EI/ ���/!�dDa�C@Nc�@��p�� 4	���EpANOGfAN1A[�ā�AIt����DCSZ���cT���bO�hO�gS?���b�hS�hNHIGN������A�(��dDYE��pTLL�q�2���*Є���T�"�$���}��Ԛ�SA������ʰ���Z�� �P1�u2�u3��q���R�`*І ���V��c��5�z��x�6��P�6�.�ST���R�0Y��`Q� _�$E_�C_��� I�n������T)ч Lo���瀖�x������_�ENS�_��t~D_ � =��h0Y���@�d�M�Ch2� ���C�LDP��TRQ�LI��D�2�FLAGZ�2�3�f���Du�f�`�LDf�P�f�O�RGjQy��(RESERV��Ŕ��Ŕ�� #�3�� �� 	O�jUA�f�SVHX0D�R	���'�RCLMC5�şן�G���'��ՠJ�/��3$DEBUGMAS��S�D�"���T�`p�E� TZ���MFRQ���� � �HRS�_RU�ځ�A<)��UFREQ� J��$``�OVER�h����v|P�AEFI��%�����r��ѣ� \ ���$U��3?����PS�p7 	�C�06�BҒ�G�9U�Н�?(����MISCi� d�q1�RQ5		TBB@�� ��aa��AX9�!	�"�EXGCES��_1ܲM��J.���9�ٵ�SC� � H���_G���,��� �2�РK���|��B@���B_�FLIC���B@QUIRExSMO��O��d�`p�ML܀M��� �
��19Э��5� T�MND�1e�/!�o2f2�x�D�#�4�INAUT(A�4R#SM� ��pNZ�b!��S^�4�f�PSTL�.� 4��LOCf�RI1P�EX���ANG�b����Zb Aե��p�x MF�%7�+��ۂ5`�e�c0��SU�P�dgf�FX�/ IGG�1 � ���ۃb!��ۃ�V ۄ��V�P���R���R������SD�w��TI�j��pb!M ���� t-�MD*��) 8��`C�L�@�H��C�DIA�D�2 W�]AC��q��C�D�3)ƚ�MOh�/� -a�CU�V������N�OPA_��.�� �/��7㉠f�	�
 ��P��>P����P��KE�RR�#-�$B�����ND2xN�ND2_TX䄏XTRA�cp`��&9�LO�0/�_&�� �i2���ܞ��RR2൜�� -��1A$� d$CALI���c%G�a�2�pRI�N�!�<$R� S�W0S� `�ABC>�D_JV ���7��_J3K
E1S�P����PEl3Pk����J`�h���OiqIM`�ŲCSKPS��� $�c�J�1ŲQ�%p�%'�_AZ#���=!ELNq�N�O�CMP�(���z0R1T��h#�1���F�1��(o`�*Z�$�SMGMP�n�JG��SCLB���SPH_�`Ű+0�#\ �=� RTER�I�`� _�`�*�aAP@G�Ų4DIS!��"23U�DF �  �=0LWB8VE�LD�IN�Z`e0_�BL�`��m4���J`]4r7�7�4N�IN� �������5QB��t�1��_̰ ��5 �2#5ٰ�4z�936FN�DHB�r ����p�$V� ���#oaa$� ����$\�m�R�����H? �$BELN 姾�!_ACCEs1 ��H`��@IRC_40���NT��/�O$PSB�7�LH0��DL��0�G3�`@�F;�I�G�C�G3�B��E�_�qPB-P3Q�ܰ��A_MG��DDPQ2��FW����C�lU�C�BaXDE�[PoPABN�GRO� EECR�q�_D�!�q������AH0$US�E_� �cP�CTER�dY�Pb@"� ��YN߰Aa`f�Z�BaM����bJPO_0�AGdINC���R�pT�ig��ENC0L��A�B��@IN7�I�B�e��$�NT]3�5NT231_@2���cLOQ0���`-�IP����fF0�� ��� ���e��C�0�fMOSIUQ����3Q��ŲPERCH  s+�2 ]w�hs ��rn���c'["e
P$2P�A�B�uL�T������e��z�vvT3RK�%ʁAY��s ��,��B;�0��n&��wbȠMOM��� �������S�G��C��R� DU�(RS_�BCKLSH_C �B����<v,�"c��݃�b�1a%CLAL�M�d��m�@�CH�K��NGLRT�Y��5�d����_�Z�1t_UM��l�Cૣ^Q�!����LMTh_L��V#��j�E��Ð�����E���H`}���r��xPCnq¡xH���TUl�CMqCv^PbWCN_�1Nuc��SFtA�yVb�g�!8��B��n<�CATs�SHZ� �bT�f]����f��A��	� QPPAs�gb_	Pr�V�_�� 3�Qp0�C�U�F�JG>�X��I�K0OGV�2TORQU�P�/sL��P`��Gr1�P��_W�� ,��!QAٴBCصHCصUI�I�IHCF$�`˱�-��ZPVC�@0����N�1T�RPh�$!Z�JRKT̙Ɩ��DB� M���MΏ�_DLBA�rGR�Vߴ��BC��HC��H�_����@�COS�p �LN��6�W� =�B@8ٵ 8�
�t�b��(���Z1�Gv��MY�?Ѳ��='���TH�ET0uNK23�HC��<C@�CB�C5B<CC� AS�'�`
�5�BC5��SBBC�S��GTS��QC�o/��'��'��q�$DUC��w���t5���5Q�q_��NE��AKS�z)!8 @��A���'����LPH����e��SW�o�b�o�q����P������V@�V5�T2@X�Vg�Vt�V��UV��V��V��V��H@�Y�_W�ܡvt�UH��H��H��H��UH��O1�O@�O�	�V�Og�Ot�O��O���O��O��O��F���"�~bՃ3�SP�BALANCE_l�ѮLEj�H_��SP�1S��b��q�PFULC�"��"q��:1�|!UT�O_>�F�T1T2B)�B2N%��B�`b$��!f� ���B}C��T��pO50�AɰINSsEG�B qREV�&� p�aDIF��91ٞ�'321�	�OB�!	��Ó�2���`0�~��LCHWAR�R�7BAB%���$MECH+���9a?1T�AX9�P�X6�#B7 � 
Y2��{A�e7ROBQpCR�B�5�M��0�CyA_A�T� � x $�WEIGH6`��$1��3X�I6a�`I9F�QjPLAG'b�qS'b� 'bBILEcODo�#p�2ST�@"�2P�!	��0 `@Ơ�1�0��0
�`yB(a�A�  2�.t�6D�EBU�3L�@<B���MMY9�E� N8��D�$D�Axq�$�@S��� � �DO_�@A�1� <�0VFL U�$(a�B&B@N�c�H�_p(`BCO� _�� %��T�`ķa��T�!~D�@TI�CK�30T1�@%NS��WPNQp1 �CQpRԀ(a!2iU!2uU�@_PROMP6cE�? $IR��&apL��R�p�RMAI��haa8b�U_@�S�� B�:`R��COD�[CFU.`�6ID_�ppe� �R�G_SwUFF
� C4a�QdRDOlW� mU @lVGRC!2Id �SUd!2`e!2le��Id��De@��0H� _F�IZA9�cORDf&A �0�B36���b&a�@$ZDT�e 	�CA�E��4 *�!L_NA�QWPriUDEF_I)xr�V5tuU-BhV�7DhVasuUou�VIS������A��hT�suS�3t���D4l���7BDP5 ���t[CD��O�>�BLOCKE�Cc�i_{_�W�qIbC`UM HerIdasIdouId�r UbK�TeDsUdtUb5F ���q`c,0B�`er`e@as`c���EhPP�  �t,P�q��@W*�)�� �	  �TE|��D� A�LOMB_C�^�0��2VIS!�ITY��2AS�O'CA_FcRI2#��� SI�q����RTP��_P��3tC�2W��W������r��_��jaEAS�3�jbd������p�R��4ꭙ5��6�3ORM�ULA_I��}G	w� h �N�7�ECOEFF_AO;Q� ��;Qr�G�2�3S�0�BCA �O��CCAGR�� � � $ �u"�BX+PTM�� �ARX(�%��CER� T	��t�`�  +"LLtkd�pS�_SV�t&w�$L��`���v��`� ��SETU�sMEA�P(`F���0CA�b�0� � ���0 �@o�� Q2��q�rWP�q��tբܑub��Q�p�q�p+���� ��PREC�a���MSK_���� P�11_USER^!�"}�08��}�^!VEL"�}��0��!1I�`J ��MTQCFGs��O  YP� OG2�NORE�0P����0��� 4 pݳB7�2H1XYZ�c�J!o yCH0 ��_ERR�1� �I�Q��Pۣ@�aAi�����@BUFINDX��I�o MOR� H�0CU@�QH1����Q�a���"�a${0��~q�@�;���G� � $SIj����P�!Ɓ�VO����0OB�JE���ADJU�B�� �AY�p5��D.�OU�`Վ�'a.�b=��T� ]�8��\��BDIRa�i�p� ��"�0DYN�$����T6 �R��,P�&@��OPWOR��� �,�@S�YSBU �SO!P��cҎ���U��� 1P ����PA���X�C2�OP^`U�!���!XB�AI�IM�AGS��0U�7BIM��o�IN��@�n�?RGOVRD��	���K�PM�m�0� ߀(�s��H2L�B=з >�PMC_E�`cъ�ANM��A�B1n�B 
���SL��t�� ��0OVSuL�&S�DEX�qD}p/2G2� ��_�� G�`��G�`Qfa�B�C�0p�%�c^��_ZER����s�� @вb5MO`RI��s0
�`�P�	��qPL����  $FRkEE��E���f�T�!�Ls����TD0�;@ATUS㰤AC#_T��r�UB�_�H��s�A4�`t��C D�AI�2RL���a2S�an S���XE@Y������ ��0XUP��p�qP!X�PF�D3�����PG�Ÿ��$SUBGb5��G��JMPWAIT8�V_%LOW�BQ��@CVF�QZPG2bb!Rz���U3CC� �R��MR�'IGNR�_PL�DBTB2;@P�qH1BW�P�$2��UP�%IG0�P=IG3TNLN�&2�R�����N�P)P�EED�8HADCOW;@�����E7pS4F1!4pSPDs�� L�0AV�5ps0�3UN�0"+0!R��LY�`� Q�e�P��v1�G�!$��M�P�@L+�NPA�T�2xD���PIP%w0���ARSIZ�T��c|q��Om`�h�ATT����"\�B$�MEM0�B�A>C�3UX��rBL`�ļ $��~�SWITCHZ"Z�AW��AS�8��CLLBv1��_ $BAZ�D�s�BAM� ���I���@J50����B6|�F�A_KNOW�34R��U!�AD�H۠�~0D��5YPAYL#OA鱱�SS_s�\WT��\WZYSL��A��mpLCL_�� !���R�A���T���VF�YCK��Z��T��I�XRM��W_Ғ�TB���J)a_�J�Q����AND�^�9�8d�R�Qw��P�L�@AL_ �@�@~0���A��k�C"�uDXSE!��J3M`�af� T��PDC�K��r�COŰ_�ALPHqc�cBE0��W�qo�l �Т�!>�� � �40R_WD_1YZ2�TDŰAR�4x!uEv0s��TIA4_y5_y6"�MOM��ks�sxsh�s�s��Bv ADksp�vxs�v�sPUB��R�t�uxs�u�r�B�p��� L$PI�1s��^W.��TxY.�I:�IH�IV��<p}Q7��!�� !���b�ӆ��73HIG�C73w%p4Іp4w% � z�І�߈�!!w%SAMP���B��ЇC�w%�@>c  5�q���7 �Ҁ� �� p0"p��0p������hp0���	���INќ� &�ؘ��ϔw"ښ���:�GAMMƕS|[%�$GET��o��D�d��
ϡI�B��2I0�$HIB�_��sЩү�E��b��A��٠ʦLW�� ���٩�ʦ�b��0:caC�%CHK��� 	��nI_%����� \bxΑ�����s���v|���c �$�h� 1���I� RCH_D��'� �$)�LE�������h�ذ�0MSWFL��$M�`SCR
(75_����3��dƧ����kp��x�p0�ĴDSVv1�P��v�K�x��	���S_SA�AX�����NO�`C� ��d����d_v_\��J�:ۂ�+R��w�0sD <�4���40��zʴ�ʈ ��چ�1����ՕәS� ��@M�� 7� ��YL,�a������-���-�� ��b��9�az�K����W�{����py�Ȳ�M� ��P��`a��$ 7��"�M���� � $����$W���ANG ]�Q���d���d���d��d� נNP���C���ϐX�0O�cΑZpq��� �� �<�OM��"��1�C�8U�g�bpCON��0�1PL�a_�B� |�a�����y7xs7 �s��dzdO~z�A��(�4��ǲ@�P�P A�PMON_�QUG� � 8��0QCOU��ǀQ�TH� HO&�� H�YSD@ES�B� U�E� ��@O5$� � �@P�৥��RU)NZY��@O��� � POP+�%���>2ROGRA��x@�:�2�Ov+ITx�xINFO���� �A_�8��v��OI�� (ʰSLEQ������zb�S_EDd N� � ���r�K�QjI#��EȠNU'�(AUT��%CO�PY�Q��8,���MⵡNB F+U�PRU�T� I"NF2U��B$G0�$�aP_RGADJ!�B3X_��2$�0�&~��&W�(P�(��&�73� �NH`_CY�C� �!NS�D���LGO�b��`NYQ_FREQ�rW����^1RD)L�P:BV0�!�s����CRE���c�I�FH�jNAK�%��4_G�STAT�U å�MAIL�I�S&@V��ǀLA�ST�1�a04ELE�M:1� �EaNAyB�0EASI&A ��v�n�?�B���GF�����I���U2��0�� �|BAB�C	PRS�LV	A�Fa�Ię��qU����JP�'c�FRMS_TR vCΑ��Ci����Af�D E��& �	SB 2�   �V��9V(b8WR��`�RNTdW&�
�DO�P0�W}��04PR �;0=��GRID}�oBARS��TY'C;	� OTO�p!W� _�4!� ��R�TOo�74� �s |� PORX�c�	bSRV�0),(d fDI��T!pAa Td��^g��^g4\i[��^g6\i7\i8@bM��PFj�:1�$VALU�C��9D�7@F65�� !!"E��l�S�1��F_@AN���b�1R |c17ATOTALH�,�qCsPWK3I�QYtREGENWzlr��X�H@c5v� T1R�C�Wq_S���wlp\CV�!���u���1GRE�3�P�6B+�.  sV_H�PDA8���p�S_Y�i��o6SV�AR��2�� �"IG_SE��3�p b�5_/�tC=_�V$CMP���KDE�M���Ie��Z��^���bENH�ANC�� p�&Q$E�2���IN�T?`iq��F%�M�ASK=��@OVR�P� �P��1Α�Wp!;�T� 4� �_XF�{�V�PSL9GV�:1� @K�� p5a���ApJpSh��4��U>�!����sTEa��`���`��U�Jd���3IL�_M~4���p� T�Q� ����@-�\�V�4�CB�P{�4AL�M�c�V1b�V1p�2��2p�3�3p�4�4p����p:����p���j�|�IN�VIAB��<�)���0�2,�U28�3,�38�4,�!48� hR�S��� ��T $MC�_F�  ���LP����ׅ7pM8�I׃���S ( ��n��KEEP_HNA�DD��!ﴙ@��C��0��Q��?��O��| ���p�܇.�REM'��IqPbL�c�h�U�4e��HPWD  ��SBM��PCOLLAB��p��5q�2�IT50`�w"{NO��FCAL�ܔ��� ,��FL|�A$SYN����M� Cq��XpU_P_DLY!��DELA?�Jq�2Y� AD��	��Q�SKIP�� �4`-O;�NT�]�i�P_-V��^U� *����q���q��u`�� �`�ڏ`�ڜ`�ک`����`��9�!�J2R�0� �L�EX�@T X3N�7AN� �N�}� RDC���� ���Rz�TOR� ���R�1�����;TRGEA�rh@�㎉RFLG�^�5�E9R���SPC�1�UM_N��2TH�2N�Q�A� ?1� �A��Q>62 � DKш<��@2_PC3]��S���1_0L10_�C}2� 2��� �� $b� ��� 	ViR����0�� �\Ub����mrj���C1��=���ID� Gy�XUVL�1a�1n��� 10c�_DS����M01��F�11!� l������#C��AT E��$�Q���f���;T�3�HOMME� �h2n�t������3n��'9�K ��i4n�n������5n���/!/3/E/,0f6n�h/z/�/X�/�/�/ e7n���/�/	??-??? +�f8n�b?t? �?�?�?�?�5S���!�  �Ag�p�����c�Ed� aTC�tD:vtCIO�ҔII@f�O��_OAP�E�C4r��e�R� {WE�� ^@��l���4t ���B$DSB��G#NA��3s:�C��`�;�RS232zE� ����5���I�CEUS=sSPE|(��aPARIT ��2qOPB���bFLOWO�TR9@?rt��UX�CUuP���aU�XT��a�ERF�ACZTT�U�`�}�SCHa� t�఩�_`Py���$L ��pOM8���A��8�𥀯�UPDư��f�qPTU@��EX��8#hc�EFA8����pBSP�P�a��|�`�7$USA�X��9��EX�PI��$(`�pY�eR_$�q�`mQ�fWR�OI�D���f��FFRI�END��L�$U�FRAMc�pTO;OLvMYH��r�LENGTH_V�TE�dI�;s��$Z pJxUFIN�V_^ ��_ARGuI%���ITI��bBwX�Sw�vG2�gG1�aꀎc�r�w�_r�O_XP��L�+q4���N�Sc��Cp�Pr�q��G���Rǁ󐒧�XQ؂� �h�U���U�Ѻ����P�Ud�X m`E[_MG`CT�cH���h���U�dScG�W$�`ć��لD]и@KȅJӂй������{$-� 2��H�an �i1�h�`2�k2=�3�k3�j-��� �iK���F�`l��`x��|�NtV�uV��Pq�(,��r�P����V� ��#���R��pr#�.���E9�<�Os)Eg$A��T�PRh��U�k�ǓS��P��8�"Sb;Q� ! ��D��"��K��"����S`�p�p��
�$�$C��S����i��9�9� ؠ�VERSI�`����i��I�#PP��AAVM�_�a2 �� 0  G�5�V�b�S�.�� ��	������9� �����ζ����ϧ��R�d��l�0�BS^ r1��� < @ϱ����������� /�A�S�e�w߉ߛ߭� ����������+�=� O�a�s������� ������'�9�K�]� o��������������� ��#5GYk}`����|�CC`�XLM�@��n��  d�IN�����qEX?��D2_`=� ����0�IOCipq ��PZXQ��{�{IO'PV 1=�P $-��ұ�!�� �?��� �� //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5GYk}� �������� 1�C�U�g�y������� ��ӏ���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�[�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ������� LARMRECOV I���LMDG K����?_IF �� �p߂ߔߦߴ�^����������, 
 �G����m������$_������ �2�D�V�h��NGTOL  I� 	 A   ������ PPINFoO %� $�������   1�I
�8r\� ������ &W�p�Rdv�� �����//*/�x�PPLICAT�ION ?�����LR Handl�ingTool �y" 
V9.1�0P/25��5'?
88340z#�*sF0�!�/131y#��,�/�"7DF1x� 5,y#None5+�FRA5/ �6�-B&_ACT7IVE��  [#���  X3UTOM�ODb0)��U5CHGAPONL�?� �3OUPLE�D 1M�� ��0�?�?�?O;CUR�EQ 1	M�  UTILL	XO�iE_ ~D��B�m%MDH�6E�2cJHTTHSKYwO��D\CO UO_�O7O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_oo#o5oGo Yoko}o�o�o�o�o�o �o1CUg y������� 	��-�?�Q�c�u��� ��󏽏Ϗ����� )�;�M�_�q������ ��˟ݟ����%�7� I�[�m����믵�ǯ ٯ�����!�3�E�W� i�{���翱�ÿտ� ����/�A�S�e�w� ���ϭϿ�������� �+�=�O�a�s߅��� �߻���������'�09�K�CETO��d?�X2DO_CLE�AN�?V4��NM ; �� O*��<�N�`�r�NDSP�DRYR��U5HI�0�@����� &8J\n����R8MAXI ��|�~A�7�X���!�2�!>X2PLUGG�0��\�3t5PRC��B�E����.O3�����SEGF�0K z������/p/&/^�LAP�� ��Cz/�/�/�/�/�/ �/�/
??.?@?R?�3TOTAL��3_USENU��;� ��?~B@RGD�ISPMMC�2�AC��@@���4�O�����3_S�TRING 1
~�;
�M�0�ST:
)A_ITwEM13F  nT= OOaOsO�O�O�O�O�O �O�O__'_9_K_]_�o_�_�_�_I/�O SIGNAL�-ETryou�t Mode4E�Inp�PSimu�lated8AO�ut�\OVE�RR�� = 10�07BIn cy�cl�U8APro?g Aborc8A��TStatus�6C	Heartb�eat2GMH �Faulug~cAler�i�_�o�o�o�o��o $6H ��/K��AOK�� ������)�;� M�_�q���������ˏݏ_WOR�/K� ��=�O�a�s����� ����͟ߟ���'��9�K�]�o�����PO-Kia��-���ܯ�  ��$�6�H�Z�l�~� ������ƿؿ����8 �2ϴ�DEV��]� ЯJτϖϨϺ����� ����&�8�J�\�n���ߒߤ߶�����PALTu}�-���)� ;�M�_�q����� ��������%�7�I�8[�m���GRI� /K ���������� '9K]o��� ��������0Ru}I��#q�� �����//%/ 7/I/[/m//�/�/�/7PREG�� a �/?'?9?K?]?o?�? �?�?�?�?�?�?�?O�#O5OGOYO�]�$A�RG_�D ?	�����A��  	]$�V	[�H]�G���W�I�@SBN_?CONFIG�P�K��Q�RQ�ACI�I_SAVE  ��TQS�@TCE�LLSETUP ��J%  OM�E_IO�]�\%MOV_HVPi_o_�REPL�_�JUT_OBACKAQ�I�QFRA:\�+ �_�&P�'`T`�'h�� k
P �18/02/09� 11:06:04�&�H�-{o�o�o�o�\���o%7I[�&��o�� ����n��+� =�O�a�s�������� ͏ߏ�|��'�9�K�p]�o���X�  �Q�_�S_\ATBCKCTL.TM�����ҟ�����[IN�I�AeV�SMESSAG!P/�Q�@�SQD�ODE_D([P$VUb�O_�q���SPAUS͠ !���K , 	���@�Eѯߧ,		ɯ��'��#� ]�G���k�������ۿ�ſ�ͤ���TSK�  ��o��PUgPDTh�-�d~��~�XWZD_ENqB-��J��STA,���A~ŎAXIS�@U�NT 2�EQ�P� 	 �sR ��k�R"0`� Q�H�Ƹ�*��/d��U�+�>�)� v��� g�� 6�_0X �� 5�!,ߍ�Pߊ�\����METK24��-S P��@h��
@K�k@�*��7���?�I�$@7|��>&�I>.�=���f5RI$<���>&+���S�CRDCFG 1��E�Q �)UR�߆��������o�*Q%Ys�0� B�T�f�x������� ������,�����G�QGR��r���k֣�NA�P�K	��Th_ED+�1�V�� 
 �%=-��EDT-Y�Zh�M�1c���(�R��*�B�otV(��)�u2~�[ \���o�Q�/Yk/�w3J/��/ ��s/�/%/7/�/[/w4?�/c?�/�??@�?�/?�?'?w5�? R?/Ov?�OvO�?�?eO�?w6�OO�OBO ��OB_�O�O1_�Ow7z_�O�__��_o U_g_�_�_w8Fo��o��oo�o!o3o�oWow9�o_�o��;��o�o�#wCR}�_*�<��] �p���_��k � ?NO_DELw��GE_UNUSE�u�IGALLO�W 1�	  � (*SYS�TEM*��	$SERV_GR���*���REG3�$8U���*�NUMX�}��k�PMUր���LAY�С�?PMPAL,����CYC1o�l�˝x�����ULSU��0l�̒��5�L�?��BOXORI\�C�UR_,�k�PM�CNV��,�1�0����T4DLI���%�G�	*PRO�GRA2�PG�_MI�����AL(¥����B�*��$FLUI_R�ESUЗX�b�����������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ����������H�k LA�L_OUT ��T�WD_AB�ORѐ��jO�IT�R_RTN  �st��O�NONS�TO� z� b�CE_RIA_I���z������F?CFG �
���s}��_PA9�G�P 1�����Q>�P�b�!�C��p����z�C�Ce ��(��C8��e@��H�� CX��U`��h��p��x}�U������������	su?����HE��ONFI���Y�3G_Pr�1�� ��ă�} �������3�KPAUSI�1`�� ���C` 1oU���� ���/5//Y/k/�Q/�/Mo�NFOw 1`�� � 	-��/�p�� ��	�@���>�"��vm��´�B���������/�C�Q�Ch@C3����ux�B����1�C�,B���Ã�I��䮵9lfw�480��O����sw��COLLECT_���&A���~7�EN z���2W1N[DE�3�7e����1234567890�7~rD����?�6ss
 ���q)9O^OD�8OJO�OE� |O�O�O�O�O�O/_�O __w_B_T_f_�_�_ �_�_o�_�_�_Ooo ,o>o�oboto�o�o�o��6B�2�; |�=�2IO  �9 �1yxy�as��/w�TR�2!}�� bJy
�o�~> ">}x�z���9_MORr�#
� �Up�C(�n/X��!X�p�^��������ʋ1� �q$J?�,C?,,��BUpK�TqJr��P[2	&�?"�+�a�s������
R���t7���u��y���5���s� ���9PDB/�(�7��dcpmid�bg�]�v o�:���nD�pI���m�  ��nG�毱���ï��.�����mg�x�C�Ůf�g����-ſ�`ud�1:���z'�DE�F 'y(Is)���c�buf.t�xt�g��%�_M%C8�)7�!sd�ōÂ7�*��������|�C�z  B3A� C����B��0C�CI<g_6�C�C��-E���D]qeD�J�0?���D�I߁Df���-F���FR��F@���Cܤ�F@?��F[�U|ɰ����,|��t7A�UpH UpH ޒH ��t
��� ќ�@ Da  D��  E	� D��@ ��;�| F�p F"� G�=�fF��G�'i�-G>��Gg� GK  �H�<=H�&�HyMc��  �>�33  `C�/��n)���5Y�T娂��A�|�=L��<#� �Vq�����ξ��RSMOFST %8ʝ/�&�P_T1��DE ;-3����q��Tq;������??���<�;��EST2�+8�PRb�2.a?����C4��%�|��Up���������C��B���C�����H�Up:d�� ���T_2�PROOG ���%x��V$INUSER�  �5($KEY_TBL  ��"�	
��� !"#$%&�'()*+,-.�/�7:;<=>?�@ABC2�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������0��͓���������������������������������耇�������������������s��q* LCKtx��&t STAT����_AUTO_D�O�6���IND��4�}1R���T927/�STO@/� TRL, LET�E�7~*_SCR�EEN ?�_kcsc�2Uo �MMENU 1/.� <ED? [�/?J?ճ'?M?�? ]?o?�?�?�?�?�?�? O:OO#OpOGOYO�O }O�O�O�O�O�O$_�O _Z_1_C_i_�_y_�_ �_�_�_o�_�_oVo -o?o�ocouo�o�o�o �o
�o�o@)v M_������ �*���9�r�I�[� �����ޏ��Ǐ�&� ���\�3�E���i�{����ڟ��ß�Ϲ�#_?MANUALs/�!�DBCO RIG��'�/�_ERRL&2 0��a�N���쵯ǯ P�NUM�LI;�Z!����
�P�PXWORK 11����'�9�K��]�o��DBTB_��! 2��ç�����DB_AW�AYX�a�GCP� ��=E�ö_AL;��òT�Yr �%��I�_r� 13#� , 
�T��B�,ω�_M I��Ѽ�@����ONTIM6�'��������
�$�MOTNE�N��z$�RECO�RD 19�� y��ψ�G�O�O� =߈�Ҳ{ߍߟ߱�H� ����O��s�(�:�L� ���߂��ߦ������ �� ���$���H���l� ~��������5���Y�  2D��h��� ������U
y �Rdv��� �?�//*/� N/9/G/�/��/�/�/ ;/�/�/q/&?�/J?\? n??}?�??�?7?�? �?O�?�?FO�?jO�? �O�O�O�O_O�OWO_�{O0_B_T_f_�OòTOLERENCдsB��ްL��P��CSS_CNST_CY 2:����	i_���_�_�_o o'o9oKoaooo�o�o �o�o�o�o�o�o#��TDEVICE ;2;�[ ��v u���������*��ϭSHNDG�D <�[�Cz||{�TLS 2=]}<�����Џ�����>��RPARAM >0� |��}��SLAVE ?�]�I�_CFG �@J�*�dMC�:\�PL%04dO.CSV)��cџl�RA ��CH��o�o�*��F��w�*�6�c�s�a�`��JPѓ�|頪��r�_CRC_OUT A]}��.��_NOCOD~�B�0���SGN �C&��&j���20-APR-�21 23:42��*�09-F�EB-18 11�:06��v LIX�v�r�*�s��Iu5�M���Þ���������VERSIO�N -�V�4.2.10��E�FLOGIC 1�D�[ 	���+�ɘ�!��PROG_ENB�e�A�WULS�� d��_ACCLIM�Ư������W?RSTJNT���*��MOJ�����INIT E�Z�&�*� ��OPT�y� ?	����
 	R575*�V+�740�61�71�)5�[�1U�21ԋ�����TO  �݉����V��DE�X��d��Hp��P�ATH ۦ��A�\��9�K�[HC�P_CLNTID� ?Ѷ�� �"S��QIAG_�GRP 2J��� Q 	 �@K�@G��?���?l��>�������Q ����ᴝP)���?�b�?PT�i��^?�Vm?S�ݘ��f40�3 678901�2345{������� ��s��@n�ȴ@i�#@d��/@_�w@Z�~�@U/@O��@I��@Dc(����@����p����PA�P,�P�B4��jp���ط�
��1��-���@)hs@$���@ bN@���@����@�D@+�ʀ��������	 ��R���@N@I��@D�@>��y@9��@4�� .v�@(��@"�\Pbt���L�@Gl��@BJ@<z��@6��0�`@�*� $N�@��� $�=q@����F@|�@�33@�R@�-?���?�?�`?�+hz�����Y"J�-@&�@N����!?�?� ��// */</�-�/?�/&? 8?�/?Z?�?^?�?�? @?R?�?�?O�?4OFO �?VO����9�QH�i @��V�AY����?�z��A���5AF�A4���@��L4R��A��@�p� R��Q�R-PP��@ِ� ��Ah��=H��9=Ƨ�=��^5=�>P���>���=��,d_�,P� �z��C��<(�U\�� 4����_����A@��?��pO�_ xM�_o0o�ȡT<ofo� ovo�o~o�o�o|I>���y�b�R=���=��zq����G�G���� � ��!�!�NUt@��T��V��uB��� B�B��B%���H����~'���u��8�q�q6|�\�&�P��g���)PB3pB�5B A�@�"����m���<��  �5�-T�6��LT��o5����5���E����C�/d�C?O�ChA��l�@��r�ݏȏ��x��"�����C3����u�lB���?H��q�쏕��������ݟȟ ����澺�Ƚ��ܷ�=��<��SxM�=����CT_CONFI�G K�m��eg7Ų�STB_F_TTS��
Yɠ��Ȱ��������M�AU��N�N�MSW�_CF\�L��  ���OCVIEWf��M��ᄀ�� A�S�e�w�������/� Ŀֿ����ϭ�B� T�f�xϊϜ�+����� ������,߻�P�b� t߆ߘߪ�9������� ��(��L�^�p�� ����G����� �� $�6���Z�l�~�����,��D�RC�N(E��!P�����!E4�iX���SBL_�FAULT O�����GPMSK����P�TDIAG� P`��qo���o�UD1:� 6789012345t�n���P*�Sew��� ����//+/=/�O/a/s/2���R
�B�/J�TRECP�
?)�+A >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO�^O�/�/�/�O�UM�P_OPTION����ATR袒��	��EPME���OY�_TEMP  _È�3B�5P9��TUNI͠���5QܦYN_BRK� Q��EDI�TOR�A�A_�R_~� ENT 1R���  ,&Z�AD15 ADR�A͠�_iH&ST�UDKW�_�_&�-BCKEDT-8	o�^�R4  %o7oR�R3Oo�o�S2{o¸o�S���o�M&STYLE1�o�bo&PROG_��o<&}bs��P�t���� ���/�A�(�e�L� �����������ʏ܏�� ��PMGDI_�ST�Q�F5Q}UNCr;�1��� �dO(��v��N
�Nd�Oݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W��En��� ������ʑ��ؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@ߺ�g�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�_� i�{������������� ��/ASew ������� +=W�Es�� ������//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?O ak?}?�?E?��?�? �?�?OO1OCOUOgO yO�O�O�O�O�O�O�O 	__-_G?Y?c_u_�_ �_�?�_�_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o%7 Q_[m��_�� ����!�3�E�W� i�{�������ÏՏ� ����/�IS�e�w� �������џ���� �+�=�O�a�s����� ����ͯ߯���'� A�3�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������9�K�U�g� yߋߥ����������� 	��-�?�Q�c�u�� ������������ ��C�M�_�q����ߧ� ��������%7 I[m���� ���!;�EW i{������� �////A/S/e/w/ �/�/�/�/�/�/�/? ?3!?O?a?s?��? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_+?=?G_ Y_k_!_�?�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	#_5_?Qcu�_ �������� )�;�M�_�q������� ��ˏݏ���-7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ���%�/�A�S�e�� q�������ѿ���� �+�=�O�a�sυϗ� �ϻ���������� 9�K�]�w����ߥ߷� ���������#�5�G� Y�k�}�������� �����'�1�C�U�g� �ߋ������������� 	-?Qcu� ������m�� );M_y���� ����//%/7/ I/[/m//�/�/�/�/ �/�/�/!?3?E?W? q{?�?�?�?�?�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O? �O+_=_O_i?__�_�_ �_�_�_�_�_oo'o 9oKo]ooo�o�o�o�o �o�o�o__#5G �os_}����� ����1�C�U�g� y���������ӏ��o �-�?�Q�ku��� ������ϟ���� )�;�M�_�q������� ��˯ݯ�	��%�7� I�c�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ���/�A�[�M�w� �ߛ߭߿�������� �+�=�O�a�s��� ������������'� 9�S�e�o��������� ��������#5G Yk}����� ���1C]�g y������� 	//-/?/Q/c/u/�/ �/�/�/�/I�?? )?;?U_?q?�?�?�? �?�?�?�?OO%O7O IO[OmOO�O�O�O�O �O�/�O_!_3_M?W_ i_{_�_�_�_�_�_�_ �_oo/oAoSoeowo �o�o�o�o�o�O�o +E_;as�� �������'� 9�K�]�o����������ɏ�o �$ENE�TMODE 1T�Fu� + �`�`�e��"��RROR_P�ROG %��%��fe�r�@�TABL/E  ��P���ß՟�@�SEV_�NUM �  ��	��@�_�AUTO_ENB�  ,��=�_N�O� U��!���  *�]��J]��]��]��+\��v�����6�FLTR"�4�HIS��a��/�_ALM 1V.�� ��d]��`+��6�H�Z�l�~�䐿��_��<�  ���[�"�պ�TC�P_VER !���!]���$EXTLOG_REQ֦s�-�'�SIZ0Ϯ"�STKM�K���$�TOL  ��aDzޢ�A "�_BWD������ض�'���DI�� WFu�� ��a��STEP�����>��OP_DOo����FDR_GRP s1X����d 	п�m�"�^�n&����c?���$,MT� ��$ ������^ӳ���^�B��I�B�ĂB���BcGA����A�R1���A��3B\�B����AIG�As� A�������:�%�^�I��m��� � @� �As��Y>(�����`
? E�� 	�����}+�������p?�*�c���@  ��@�33@�������@���L�����^�F@ ������������L�FZ�!D�`�D��� BT��@��=���?�  M���6���u���5�Zf5�ES������'R��� ���`��X����2��x�FEATURE� YFu��&��LR Han�dlingToo�l ��bEn�glish Di�ctionary��4D St� a�rd��Anal?og I/O#,�gle Shif�t?uto So�ftware U�pdatedma�tic Back�up�	�ground Edit� ~�Camera:�F>Common� calib U�I��n��Mo�nitor�tr~� ReliabS��DHCP��
D�ata Acqu�is�%)iagn�os�7?+ocu�ment Vie�we"''ual �Check Sa�fety��ha�nced��
�%s� Fr��xt.� DIO �fi�u$�'end� ErEr Lt"	=�'s9�r5�  ���
FCTN Menu� �v##[7TP In�J0facq5�Gi�gE�>�5�p Mask Exc� �g�'HT�0Pro�xy Sv�$�6i�gh-Spe� S�ki��6m � mm�unic�onsHurh0J0:/;�2�connect �2:Hncr�0st#ru8Ja@e�!� �Jt%�KAREL Cmd. L�0�ua�8�CRun-;Ti� Env�HK0�el +�s�S�/W�Licen�se�#�,0Boo�k(System�)�
MACROs�,�2/Offse�ZUH� w8/"PMR �s.M}M@!�l�,MechSt�op�1tQ@Y"Ui2V�Vx� 7�L^�odTwitch��_aSh!.BV�[OpctmoaS�0fi�^�aVg0GUulti�-T�0��	PCMO funkG�ia�P�tiz~h�goV$R�egiPr@�fr�i� F�k�f8Num Sel�U�i�  Adju@�n q<V1}tatu�aI��*�RDM Ro�botscov�e�ueav`� F�req AnlyNGRem�P�!n|�u�rServo� ��P�SNPX b��B[SN�0Clix�!�WLibrD(��  �T:��vo�@=th0ssag~e��� l5Q&�/I|�=��MILIB��~��P Firmu:��Ph3Acc���TPTX4/��el�n5PǏ���1U��o�rquTimul�a!�E�u�PPa��A���!!c&�0e3v.��mri� ��USR EVN�Tğ֐nexcept� �pn�#ѕ�(@VC�rBB�X�VU 6��G�:�A�S��SC�y�SGE쎯��UI&Web Pl`vǮ�q0O���0�$�!?6ZDT �ApplD�
iP�0a!�:� Gri=d�qplay=����W�R-�.��h!�N��B^P}200i<V4+scii�1r�Load� �Up�l���f@I�Pat�V�ycS�B�`��� \6RL��� ۩�5�MI Dev�@ �(�qR�f�?�gss�wo!�_64M?B DRAMM����FRO�Ͼell�:�sh��#�c�.k �rp��5�tyBSs
r7̬r'`.?+`�p�!"=-o� 2�=a5port�.�p4�r q�-T1 �{x]P��No m�p�c$筴OL��S�up��Fa�hOPCg-UA�l�T �2�eϓ�S0�0cro�a|�s:����~���uWest�uS��e2'texV��up�1�#Ɣ�PP�00�oVi�rt�!�sR�std�pnÛ�� SWI�MEST f F	0����������� ������ MD Vpz����� �
I@Rl v������/ //E/</N/h/r/�/ �/�/�/�/�/??? A?8?J?d?n?�?�?�? �?�?�?O�?O=O4O FO`OjO�O�O�O�O�O �O_�O_9_0_B_\_ f_�_�_�_�_�_�_�_ �_o5o,o>oXobo�o �o�o�o�o�o�o�o 1(:T^��� ����� �-�$� 6�P�Z���~������� Ə����)� �2�L� V���z�������� ���%��.�H�R�� v������������� !��*�D�N�{�r��� �������޿��� &�@�J�w�nπϭϤ� ����������"�<� F�s�j�|ߩߠ߲��� �������8�B�o� f�x���������� ���4�>�k�b�t� ������������ 0:g^p�� ����	 , 6cZl���� ��/�/(/2/_/ V/h/�/�/�/�/�/�/ ?�/
?$?.?[?R?d? �?�?�?�?�?�?�?�? O O*OWONO`O�O�O �O�O�O�O�O�O__ &_S_J_\_�_�_�_�_ �_�_�_�_�_o"oOo FoXo�o|o�o�o�o�o �o�o�oKBT �x������ ���G�>�P�}�t� ������������� �C�:�L�y�p����� �����ܟ���?� 6�H�u�l�~������� �د���;�2�D� q�h�z�������ݿԿ � �
�7�.�@�m�d� vϣϚϬ��������� �3�*�<�i�`�rߟ� �ߨ����������/� &�8�e�\�n���� ����������+�"�4� a�X�j����������� ������'0]T f������� �#,YPb� �������/ /(/U/L/^/�/�/�/ �/�/�/�/�/??$? Q?H?Z?�?~?�?�?�? �?�?�?OO OMODO VO�OzO�O�O�O�O�O �O_
__I_@_R__ v_�_�_�_�_�_�_o ooEo<oNo{oro�o �o�o�o�o�o A8Jwn��� ������=�4��F�s�j�|�����̍�  H55�1���2�R78�2�50�J61�4�ATUP�5�45�6�VCA�M�CUIF�2�8H�NRE�52�;�R63�SCH��DOCV��CS]U�869�0��EIOCl�4��R{69;�ESET$�v:�J7:�R68��MASK�PRXuYT�7�OCO�3$������37�J�6
�53��He�L{CH�OPLG$��0O�MHCR �SMATk�MCS�#�0��55�MD�SW�B�OPB�M�PRC���s�0�PCMS�5J�������s�51/�51{�0n/�PRS�697��FRDG�FREQn�MCN�93��SNBAx�f�SH�LB�M
ǀ���2��HTC#�TMI�L􈳖TPA˖T7PTX<�EL۶��ⳗ8�����J95�_�TUTC�UEV��UEC�UFR�G�VCC��OǦV�IPG�CSCk�C�SGk���I�WE�B#�HTT#�R6lv���CG6�IG�oIPGS\�RCGƻDGB�H75/�Ru7�Ry�R66O��2O�R6�R55���4��5��D06:�F�CLI3�.��CMS˖0�#�ST-Y��TO7�7��t��_�ORSǦ��Mn��NOM˖OL��$���OPIs�SE�ND�L��Sy�EcTSsּ�S�CPk�wFVR˖IPNG�Gene�È6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p������	  H�551��2�
R�782�50�	J�614�	ATUP�5456�	V�CAM�	CUIFv28lNRE�
�52[R63�S{CH�	DOCV�wCSU�
869�0+EIOC�4�R69[ESE�T<ZJ7ZR6�8�
MASK�	P�RXY|7�
OC�OL,3<X 3��*J653�H��,LCH�*OPL�G<0�*MHCR��*SJ;MAT�MkCS;0[+55+�MDSW�;�+OP��+MPR�*��,0.PCM{5KX �+X0�+51K51�[L0KPRSK+6�9�*FRDkFR�EQ�
MCN�
9=3SNBA��+/SHLB�JM[���<2HTC;T�MIL��TPA�*TPTX\ZEL��JX0�8
�
J�95�TUT�*U�EVK*UEC�*U�FRkVCC+lO�k:VIPkZCSCN�ZCSG��I�	wWEB;HTT;�R6��\CG�kI�G�kIPGS�jR�CkZDG�+H75�KR7:+RYLR6�6�,2�*R6�R�55k|4�[5�{D�06+F�|CLI�<JCMS*�p;�STY[kTO�k78���ORSk:x �M�LNOM*OqL�;�0�OPI�j�SEND�
L:kS�Y�ETS�j {[C�P�FVR*IP=NkZGene�� R�d�v���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P�bt������� STD�LANG��	 '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�Z�RBT�OPTN�_�_�_�_�_DPN�oo*o<oNo `oro�o�o�o�o�o�o��oted ��>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|����������0�B�  �K�i�{�������Í�99ʅ�$FE�AT_ADD ?_	�������?  	ǈ� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O��O�DEMO �Y��    ǈ1]'_9_f_]_o_�_ �_�_�_�_�_�_�_,o #o5oboYoko�o�o�o �o�o�o�o�o(1 ^Ug����� ���$��-�Z�Q� c�������Ə��Ϗ� � ��)�V�M�_��� ������˟��� �%�R�I�[������ ����ǯ����!� N�E�W���{������� ÿݿ����J�A� Sπ�wω϶ϭϿ��� �����F�=�O�|� s߅߲ߩ߻������ ��B�9�K�x�o�� ������������ >�5�G�t�k�}����� ��������:1 Cpgy���� � �	6-?l cu������ �/2/)/;/h/_/q/ �/�/�/�/�/�/�/? .?%?7?d?[?m?�?�? �?�?�?�?�?�?*O!O 3O`OWOiO�O�O�O�O �O�O�O�O&__/_\_ S_e_�_�_�_�_�_�_ �_�_"oo+oXoOoao �o�o�o�o�o�o�o�o 'TK]�� �������� #�P�G�Y���}����� ����׏����L� C�U���y�������ܟ ӟ��	��H�?�Q� ~�u�������دϯ� ���D�;�M�z�q� ������Կ˿ݿ
�� �@�7�I�v�m�ϙ� ������������<� 3�E�r�i�{ߕߟ��� ��������8�/�A� n�e�w�������� �����4�+�=�j�a� s��������������� 0'9f]o� �������, #5bYk��� �����(//1/ ^/U/g/�/�/�/�/�/ �/�/�/$??-?Z?Q? c?}?�?�?�?�?�?�? �? OO)OVOMO_OyO �O�O�O�O�O�O�O_ _%_R_I_[_u__�_ �_�_�_�_�_oo!o NoEoWoqo{o�o�o�o �o�o�oJA Smw����� ����F�=�O�i� s�������֏͏ߏ� ��B�9�K�e�o��� ����ҟɟ۟���� >�5�G�a�k������� ίůׯ����:�1� C�]�g�������ʿ�� ӿ ���	�6�-�?�Y� cϐχϙ��Ͻ����� ���2�)�;�U�_ߌ� �ߕ��߹�������� .�%�7�Q�[���� �����������*�!� 3�M�W���{������� ��������&/I S�w����� ��"+EO| s������� //'/A/K/x/o/�/ �/�/�/�/�/�/?? #?=?G?t?k?}?�?�? �?�?�?�?OOO9O COpOgOyO�O�O�O�O �O�O_	__5_?_l_ c_u_�_�_�_�_�_�_ ooo1o;oho_oqo �o�o�o�o�o�o
 -7d[m�� �������)� 3�`�W�i�������̏ ÏՏ����%�/�\� S�e�������ȟ��џ �����!�+�X�O�a� ������į��ͯ��� ��'�T�K�]����� ������ɿ������ #�P�G�Yφ�}Ϗϼ����������  �+�=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C Ugy����� ��	-?Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O_Y  XQ/_ A_S_e_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� ����������/ ASew���� ���+=O as������ �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O@�O�O�O�O	_QPX3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝπ����������	����$FEAT_DEMOIN  ԫ�K��!�3�I�NDEX@�Oш�3�ILECOMP Z������N�.�w�SETUP2 [������  N� ��t�_AP2B�CK 1\�� � �)�����%���!����H�� ��t���'����]� ����(���L���p� �����5�����k�  ��$��1Z��~ ��C�g�� 2�Vh��� ?��u
/�./@/ �d/��/�/)/�/M/ �/�/�/?�/<?�/I? r??�?%?�?�?[?�? ?O&O�?JO�?nO�O O�O3O�OWO�O�O�O "_�OF_X_�O|__�_ �_A_�_e_�_o�_0o �_To�_ao�oo�o=o �o�oso�o,>�o b�o��'�K��o������P��� 2��*.VR�g��p*j����s0�����uQ�PC�>�pFR6:֏���;�ʋT_�_�q�� �\���B�,����vG*.FT���q	�������C�қSTM c�l�w��d�����piPend�ant Pane	l��қH�������p��3�L�ӚGIFV������l�)�;�пӚJPGڿϋ�𿭿���T�ˊJS^χ��p��u�2�%
JavaScript��޿CS��ߊ��ϵ�� %Casca�ding Sty�le Sheet�s7ߩp
ARGN?AME.DTf��|��\z�8ߚ��Ի��g���DISP* �ߔߎ���>���0�?����	PANEL15��%�����ﵯǯu�2����������o�z�3;������L�^���z�4��%�������wr�TPEINS.XML~��:\�PbCu�stom Too�lbar���PA?SSWORDC�~?FRS:\�� %Passw�ord ConfCigW��4�/�� �[U�/qֱ䘯� ��/�b_/v���/%J(�/g/y/?'2T/=?H(+?�/�/�? ��?�/U5�?o?�?O'3\?EOH(3O�?O �O���O�?]E�OwO�O_'4dOM_H(;_�O _�_�_�OeU�__ �_&o�Jo�no�� �o3o�oWo�o�o�o" �oFX�o|�� A�e���0�� T��M������=�ҏ �s����,�>�͏b� 񏆟�'���K���o� ٟ���:�ɟ^�p��� ��#���ʯY��}�� ����H�ׯl���e��� 1�ƿU������ ϯ� D�V��z�	Ϟ�-�?� ��c��χ���.߽�R� ��v߈�߬�;����� q���*����`��� ���}��I���m�� ���8���\�n���� !���E�W���{��� 	F��j����/ �S����B ��x�+���a�,�$FIL�E_DGBCK �1\������ < ��)
SUMMA�RY.DG/�]M�D::/z/�D�iag Summ�ary{/([CONSLOGp/S/e!�/��/�!Conso?le log�/�\?TPACCN�/Y?�%A?~?�%TP �Accounti�n ?�Y@6:IP�KDMP.ZIP��?�
�?O�%�0E�xception�O�*�_\O��bQJO�_1FR DT Files�O��<f MEMCHECCKt?�/i/_1�Memory D�ata_�
l?�)	FTP�/f_��Oj_W1mme�`TBD�_�L �>I)ETHERNET�_��A�_�o�!Ether�net 0fig�ura&O�}QDCSVRF�_m__�o�Q%]` ve�rify all��o�M.cXeDIFF�ovo�o P�%�hdiff��g�A]`CHG01�o��a5��b- `y2�� &�1��gr3����� <�я`��VTRNDIAG.LS֏����.�z!Q� Ope>c� Log �!no�stic���)VDEV�DA}O�����a�VisQ�DevisceX�e�IMG��?����4�7�ʔI�mag֟c�UP�{�ESz��FR�S:\z��O@Up�dates Li�st���"�FL?EXEVENo��%�>��a� UI�F Ev�QU�?� � ,�sz)
P�SRBWLD.C	Mj��������0�PS_ROBOW�EL�_�*�HADOW4��+�D�S�Shadow �Chang�O���a��RCME�RR<�!�3���S���CFG Err{orАtailkϟ ��B��SGLIB�ϧϹ�N�:!Q� St?`_������):�Z�DU_��7���WZMDT�adn����NOTIbo�߽�R��UNotifiqc?b��t��AGXbGIGE��/�A���]�GigEZ�d��N�A��-��Q� �^������:����� p���);��_�� ��$�H�l� �7�[m��  ��V�z/!/ �E/�i/�v/�/./ �/R/�/�/�/?�/A? S?�/w??�?�?<?�? `?�?�?O+O�?OO�? sO�OO�O8O�O�OnO _�O'_9_�O]_�O�_ _�_�_F_�_j_�_o �_5o�_Yoko�_�oo �o�oTo�oxo�o C�og�o��,� P�����?�Q� �u����(���Ϗ^� 󏂏�)���M�܏q� �����6�˟ݟl�� ��%���2�[���� ����D�ٯh������ 3�¯W�i�������� @����v�Ϛ�/�A� пe����ϛ�*Ͽ�N� ���τ�ߨ�=���J� s�ߗ�&߻���\��� ���'��K���o�� ��4���X������ #���G�Y���}���� ��B���f�����1 ��U��b��>���t	�$F�ILE_FRSP�RT  ���� ����$MDONLY �1\8�  
 ��{���� ����///�S/ �w/�//�/</�/�/ r/?�/+?�/8?a?�/ �??�?�?J?�?n?O O�?9O�?]OoO�?�O "O�OFO�O�O|O_�O 5_G_�Ok_�O�_�_0_ �_T_�_�_�_o�_Co��_Poyo"VISB�CKV@e*.�VD�o�o8`FR�:\�`ION\DOATA\�o[b8`�Vision VD file�o o>Pfot^o�' ��]���(�� L��p�����5�ʏ ܏�� ���$���5�Z� �~������C�؟g� ������2���V�h�#� �����?����u�
� ��.�@�ϯd�󯈿��)���LUI_C�ONFIG ]�8�aɻ $ ��[{8 �2��D�V�h�zψ��|x ������������
ܠ� -�?�Q�c�u�߆߫� �������ߊ��)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi  ������~ /ASe��� ���h�//+/ =/O/�s/�/�/�/�/ �/d/�/??'?9?K? �/o?�?�?�?�?�?`? �?�?O#O5OGO�?kO }O�O�O�O�O\O�O�O __1_C_�Og_y_�_ �_�_�_X_�_�_	oo -o�_>ocouo�o�o�o Bo�o�o�o)�o M_q���>� ����%��I�[� m������:�Ǐُ� ���!���E�W�i�{� ����6�ß՟���� ���A�S�e�w��� � ����ѯ������+� =�O�a�s�������� Ϳ߿�Ϛ�'�9�K� ]�oρ�ϥϷ����� ���ϖ�#�5�G�Y�k� }�ߡ߳��������� ���1�C�U�g�y�	����x����$F�LUI_DATA ^�������R�ESULT 2_����� �T��/wizar�d/guided�/steps/Expert��"�4� F�X�j�|���������������Cont�inue wit�h G��ance ��1CUgy�`����� ���-����0 �������$���ps�o��� �����/#/5/ ���\/n/�/�/�/�/ �/�/�/�/?"?4?F>�$(:Jrip�X�?�?�?�?O O*O<ONO`OrO�OC/ �O�O�O�O�O__&_ 8_J_\_n_�_�_Q?c?ȭ_�?EJ�Ti�meUS/DST �_"o4oFoXojo|o�o�o�o�o�o��Enabl
.@ Rdv�����
��� �_��_�_f24or����� ����̏ޏ����&� �o�o\�n��������� ȟڟ����"�4�����)�;�M�zon 
`7�ʯܯ� ��$��6�H�Z�l�~���E�ST Ea�rn? Stand���� ��ӿ���	��-�?�`Q�c�uχ�� ���t�f�x�:���acces�?�+�=� O�a�s߅ߗߩ߻��������nect �to Network���%�7�I�[� m���������ȅ�B��Ϻ��ϊ�!���`Introd?uction��t� �������������� (�OL^p�� ����� $5�_�P*����V?Editor5� ���
//./@/R/�d/v/5 Touc�h Panel �� (recommen�P)�/�/�/ �/�/?#?5?G?Y?k?�}?�̬P�^�?���  �s/Reg `�O%O7OIO[OmOO��O�O�O�O6�EuropM�__&_8_J_ \_n_�_�_�_�_�_�_ B�z��?o�?�?��EU�_no�o �o�o�o�o�o�o�o�"��C���Ban CeX�al,ew ���������+��V�L�o	oo -o?o������Ώ��� ��(�:�L�^�p�3 ������ʟܟ� �� $�6�H�Z�l�~�:��Q�KY�k�}�����/currNp���,�>� P�b�t���������ο���14-FEB-�18 05:03 PMԿ��/�A� S�e�wωϛϭϿ���:�7�����į֯���Yea�j�|ߎ� �߲�����������>��2018(�Q� c�u���������0����)� 
���  ��f�(�:�>��Month+��� ������,>Pbt��2|�� ���� 2D Vhz9�K��S\�n�8������Day/ $/6/H/Z/l/~/�/�/8�/�/��14�/�/ 	??-???Q?c?u?�?@�?�?�?�?���pO����HouY� fOxO�O�O�O�O�O�O�O__�5$_J_\_ n_�_�_�_�_�_�_�_ �_o"o�?� Obo�$O6O��inute 'o�o�o�o�o) ;M_q�3x� �����
��.�@@�R�d�v�5o�To0��xo�o��AM��� �1�C�U�g�y����� �����)�����'� 9�K�]�o���������ɯ������Ϯ����ҏ�NetMethodϯa�s��� ������Ϳ߿����0�Not configureO� R�d�vψϚϬϾ��� ������%���� ���!���ߚ߬߾� ��������*�<�N�`�r� �ߗ����� ������'�9�K�]� o�����b�L�Xߺ� |�����);M _q����x�� �%7I[m ���������� /��3/E/W/i/{/�/ �/�/�/�/�/�/?� ?A?S?e?w?�?�?�? �?�?�?�?OO�:O �^O /�O�O�O�O�O �O�O__'_9_K_]_ o_�O�_�_�_�_�_�_ �_o#o5oGoYoko*O �oNO�orO�o�o�o 1CUgy�� ���_��	��-� ?�Q�c�u��������� |oޏ�o��oƏ;�M� _�q���������˟ݟ ����7�I�[�m� �������ǯٯ��� �Ώ0��T�f�*��� ����ÿտ����� /�A�S�e�$��ϛϭ� ����������+�=� O�a� �j�D��߸�z� ������'�9�K�]� o�����v����� ���#�5�G�Y�k�}� ������r߼ߖ���
 ��1CUgy�� �����	��- ?Qcu���� ���/�������� \/�/�/�/�/�/�/ �/??%?7?I?[? ?�?�?�?�?�?�?�? O!O3OEOWOiO(/:/ L/�Op/�O�O�O__ /_A_S_e_w_�_�_�_ l?�_�_�_oo+o=o Ooaoso�o�o�o�ozO �O�O �O'9K] o������� ��_�5�G�Y�k�}� ������ŏ׏���� �o.��oR�y����� ����ӟ���	��-� ?�Q�c�t��������� ϯ����)�;�M� _����B���f�˿ݿ ���%�7�I�[�m� ϑϣϵ�t������� �!�3�E�W�i�{ߍ� �߱�p��ߔ��߸��� /�A�S�e�w���� �����������+�=� O�a�s����������� ������$��HZ �������� �#5GY�} �������/ /1/C/U/^8�/ �/n�/�/�/	??-? ??Q?c?u?�?�?�?j �?�?�?OO)O;OMO _OqO�O�O�Of/�/�/ �O�O�/%_7_I_[_m_ _�_�_�_�_�_�_�_ �?!o3oEoWoio{o�o �o�o�o�o�o�o�O�O �O�OP_w��� ������+�=� O�os���������͏ ߏ���'�9�K�]� .@��dɟ۟� ���#�5�G�Y�k�}� ����`�ůׯ���� �1�C�U�g�y����� ��n����������-� ?�Q�c�uχϙϫϽ� �����ϲ��)�;�M� _�q߃ߕߧ߹����� �����"��F��m� ������������ �!�3�E�W�h�{��� ������������ /AS�t6�Z� ����+= Oas���h�� ��//'/9/K/]/ o/�/�/�/d�/��/ ��/#?5?G?Y?k?}? �?�?�?�?�?�?�?� O1OCOUOgOyO�O�O �O�O�O�O�O�/_�/ <_N_Ou_�_�_�_�_ �_�_�_oo)o;oMo Oqo�o�o�o�o�o�o �o%7I_R_ ,_v�b_���� �!�3�E�W�i�{��� ��^oÏՏ����� /�A�S�e�w�����Z �~ȟ��+�=� O�a�s���������ͯ ߯񯰏�'�9�K�]� o���������ɿۿ� ����П�D��k�}� �ϡϳ���������� �1�C��g�yߋߝ� ����������	��-� ?�Q��"�4ϖ�XϽ� ��������)�;�M� _�q�����T߹����� ��%7I[m ��b�t����� !3EWi{� ��������/ //A/S/e/w/�/�/�/ �/�/�/�/�?�:? �a?s?�?�?�?�?�? �?�?OO'O9OKO\? oO�O�O�O�O�O�O�O �O_#_5_G_?h_*? �_N?�_�_�_�_�_o o1oCoUogoyo�o�o \O�o�o�o�o	- ?Qcu��X_� |_��_��)�;�M� _�q���������ˏݏ o�%�7�I�[�m� �������ǟٟ럪 ��0�B��i�{��� ����ïկ����� /�A� �e�w������� ��ѿ�����+�=� ��F� �jϔ�V����� ������'�9�K�]� o߁ߓ�R��������� ���#�5�G�Y�k�}� ��NϘ�rϼ����� �1�C�U�g�y����� ����������	- ?Qcu���� ���������8�� _q������ �//%/7/��[/m/ /�/�/�/�/�/�/�/ ?!?3?E?(�? L�?�?�?�?�?OO /OAOSOeOwO�OH/�O �O�O�O�O__+_=_ O_a_s_�_�_V?h?z? �_�?oo'o9oKo]o oo�o�o�o�o�o�o�O �o#5GYk} �������_
� �_.��_U�g�y����� ����ӏ���	��-� ?�P�c�u��������� ϟ����)�;�� \����B�����˯ݯ ���%�7�I�[�m� ���P���ǿٿ��� �!�3�E�W�i�{ύ� L���p��ϔ����� /�A�S�e�w߉ߛ߭� �����ߢ���+�=� O�a�s������� ��� ���$�6���]� o��������������� ��#5��Yk} ������� 1��:��^�J� �����	//-/ ?/Q/c/u/�/F�/�/ �/�/�/??)?;?M? _?q?�?B�f�?�? �OO%O7OIO[OmO O�O�O�O�O�O�/�O _!_3_E_W_i_{_�_ �_�_�_�_�?�?�?�? ,o�?Soeowo�o�o�o �o�o�o�o+�O Oas����� ����'�9��_
o o~�@o����ɏۏ� ���#�5�G�Y�k�}� <����şן���� �1�C�U�g�y���J� \�n�Я����	��-� ?�Q�c�u��������� Ͽ�����)�;�M� _�qσϕϧϹ����� ������"��I�[�m� ߑߣߵ��������� �!�3�D�W�i�{�� ������������� /���P��t�6ߛ��� ��������+= Oas�D��� ��'9K] o�@��d����� �/#/5/G/Y/k/}/ �/�/�/�/�/��/? ?1?C?U?g?y?�?�? �?�?�?��?�O*O �/QOcOuO�O�O�O�O �O�O�O__)_�/M_ __q_�_�_�_�_�_�_ �_oo%o�?.OORo |o>O�o�o�o�o�o�o !3EWi{:_ �������� /�A�S�e�w�6o�oZo ��Ώ�o����+�=� O�a�s���������͟ ����'�9�K�]� o���������ɯ���� ���� ��G�Y�k�}� ������ſ׿���� �ޟC�U�g�yϋϝ� ����������	��-� ����r�4��߽߫� ��������)�;�M� _�q�0ϕ������� ����%�7�I�[�m� �>�P�b��������� !3EWi{� ������� /ASew��� �������/��=/ O/a/s/�/�/�/�/�/ �/�/??'?8/K?]? o?�?�?�?�?�?�?�? �?O#O�DO/hO*/ �O�O�O�O�O�O�O_ _1_C_U_g_y_8?�_ �_�_�_�_�_	oo-o ?oQocouo4O�oXO�o |O~o�o);M _q������_ ���%�7�I�[�m� �������Ǐ�o菪o ���E�W�i�{��� ����ß՟����� �A�S�e�w������� ��ѯ�����؏"� ��F�p�2�������Ϳ ߿���'�9�K�]� o�.��ϥϷ������� ���#�5�G�Y�k�*� t�N����߄������ �1�C�U�g�y��� ���������	��-� ?�Q�c�u��������� |ߎߠ߲���;M _q������ ���7I[m ������� /!/����f/(�/ �/�/�/�/�/�/?? /?A?S?e?$�?�?�? �?�?�?�?OO+O=O OOaOsO2/D/V/�Oz/ �O�O__'_9_K_]_ o_�_�_�_�_v?�_�_ �_o#o5oGoYoko}o �o�o�o�o�O�o�O
 �O1CUgy�� �����	��, ?�Q�c�u��������� Ϗ�����o8��o \���������˟ݟ ���%�7�I�[�m� ,�������ǯٯ��� �!�3�E�W�i�(��� L���p�r������ /�A�S�e�wωϛϭ� ��~�������+�=� O�a�s߅ߗߩ߻�z� �ߞ� ����9�K�]� o����������� �����5�G�Y�k�}� �������������� �����:d&�� �����	- ?Qc"����� ���//)/;/M/ _/hB�/�/x�/ �/??%?7?I?[?m? ?�?�?�?t�?�?�? O!O3OEOWOiO{O�O �O�Op/�/�/�/_�/ /_A_S_e_w_�_�_�_ �_�_�_�_o�?+o=o Ooaoso�o�o�o�o�o �o�o�O�O�OZ _������� ��#�5�G�Y�o}� ������ŏ׏���� �1�C�U�g�&8J ��nӟ���	��-� ?�Q�c�u�������j� ������)�;�M� _�q���������x�ڿ ������%�7�I�[�m� ϑϣϵ��������� � �3�E�W�i�{ߍ� �߱����������ʿ ,��P��w���� ����������+�=� O�a� ߅��������� ����'9K] �~@�d�f�� �#5GYk} ���r����/ /1/C/U/g/y/�/�/ �/n�/��/?�-? ??Q?c?u?�?�?�?�? �?�?�?O�)O;OMO _OqO�O�O�O�O�O�O �O_�/
?�/._X_? _�_�_�_�_�_�_�_ o!o3oEoWoO{o�o �o�o�o�o�o�o /AS_\_6_�� l_�����+�=� O�a�s�������ho͏ ߏ���'�9�K�]� o�������dv�� ���#�5�G�Y�k�}� ������ůׯ����� �1�C�U�g�y����� ����ӿ���	�ȟڟ �N��uχϙϫϽ� ��������)�;�M� �q߃ߕߧ߹����� ����%�7�I�[�� ,�>Ϡ�b��������� �!�3�E�W�i�{��� ��^߰������� /ASew��� l�������+= Oas����� ��/'/9/K/]/ o/�/�/�/�/�/�/�/ �/� ?�D?k?}? �?�?�?�?�?�?�?O O1OCOUO/yO�O�O �O�O�O�O�O	__-_ ?_Q_?r_4?�_X?Z_ �_�_�_oo)o;oMo _oqo�o�o�ofO�o�o �o%7I[m ��b_��_�� �o!�3�E�W�i�{��� ����ÏՏ����o� /�A�S�e�w������� ��џ������"� L��s���������ͯ ߯���'�9�K�
� o���������ɿۿ� ���#�5�G��P�*� tϞ�`���������� �1�C�U�g�yߋߝ� \���������	��-� ?�Q�c�u���X�j� |ώ�����)�;�M� _�q������������� ����%7I[m ������� ������B�i{� ������// //A/ e/w/�/�/�/ �/�/�/�/??+?=? O? 2�?V�?�? �?�?OO'O9OKO]O oO�O�OR/�O�O�O�O �O_#_5_G_Y_k_}_ �_�_`?�_�?�_�?o o1oCoUogoyo�o�o �o�o�o�o�oo- ?Qcu���� ����_��_8��_ _�q���������ˏݏ ���%�7�I�m� �������ǟٟ��� �!�3�E��f�(��� L�N�ïկ����� /�A�S�e�w�����Z� ��ѿ�����+�=� O�a�sυϗ�V���z� ���ϲ��'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� ���@��g�y����� ����������	- ?��cu���� ���);�� D��h�T���� �//%/7/I/[/m/ /�/P�/�/�/�/�/ ?!?3?E?W?i?{?�? L^p��?�OO /OAOSOeOwO�O�O�O �O�O�O�/__+_=_ O_a_s_�_�_�_�_�_ �_�_�?�?�?6o�?]o oo�o�o�o�o�o�o�o �o#5�OYk} �������� �1�C�oo&o��Jo ����ӏ���	��-� ?�Q�c�u���F���� ϟ����)�;�M� _�q�����T���x�گ ����%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ������Ϧ��ʯ ,��S�e�w߉ߛ߭� ����������+�=� ��a�s������� ������'�9���Z� �~�@�B��������� ��#5GYk} �N����� 1CUgy�J� �n����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�??)?;?M? _?q?�?�?�?�?�?�? ���
O4O�[OmO O�O�O�O�O�O�O�O _!_3_�/W_i_{_�_ �_�_�_�_�_�_oo /o�?8OO\o�oHO�o �o�o�o�o+= Oas�D_��� ����'�9�K�]� o���@oRodovo؏�c��$FMR2_G�RP 1`���� �C�4  B��p	 ��p�0��F;@ F�E��Q�F����C��L�FZ�!D�`�D��� BT��@��=�^�?�  ������6������5�Zf5�EySΑ^�A�  ����BH��\��@�/33@�� ���!�@�Q��@�g��]�Q����<�z��<�ڔ=7��<�
;;�*��<��^�8ۧ��9k'V8���8���7ג	8(��~���� �=�(�a�L����w�_CFG a��T0���ӿ�����N�O �
F�0+� 0���RM_�CHKTYP  ��p	�����R{OMF�_MINL���s��x��7�X��SSB��b��? �����u�����ϝ�TP_�DEF_OW  ��t	���IRC�OMK����$GE�NOVRD_DOrm��q*�THRm�� dG�d0�_EN�B� 0�RAV�C��c���� ��>�����v���^�����.� ��OUU��i�3�.��.�<u������,�z����sC� � D����l��$�@��B�/��1�m�\�ϑ�SMT��j���������$HOS�TC��1k���s��� MC�t�����v _ 27.0 1��  e��BTf x�
0�������	anonymous4FX@j|�r����� ����)
//./@/ R/�v/�/�/�/�i/ �/??*?<?N?� ���?�/�?��?�? OO�/�?JO\OnO�O �?�O�/�O�O�O�O_ S?�Ow?�?j_�O�?�_ �_�_�_�_+Ooo0o BoTow_�O�O�o�o�o �o�o'_9_K_]__o5 �_t�����_� ���(�K}o�op� ���������o1 3�$�gH�Z�l�~��� ���Ɵ؟����Q� �D�V�h�z���Ϗ� 󏥯���;��.�@� R�d������������ �%���*�<�N�`� ����ǯ��ۿ����� ��&�i�J�\�n߀� �ߵ�7�����������"�o���ENT 1�l���  P!\��s�  v�a� ���������
��� ���?�d�'���K��� o�����������*�� Nr5�Yk� ����8�1 n]�U�y�� ��/4/�X//|/ ?/�/c/�/�/�/�/�/�?�/B?:QUICC0O?+?=?�?a4A1�?{?�?�?a42�?��?�?>O!ROU�TER?OO-O�O!?PCJOG�OjO�!192.168.0.10h?~]3CAMPRT�O�O!�E1�@_�F�RTXO
__}_C�N�AME !P�!�ROBO�O�_S_CFG 1kP�� �A�uto-star�ted��FTP��a�Ϧ�Ao��eo wo�o�o�oF��o�o�o *o�oOas� ��r��_oo�' Io�<�N�`�r�5�� ����̏ޏ����&� 8�J�\�n�g�yϋϝ� 鏿�����"�4�F� 	�j�|�������՟W� �����0�B����� ���������ҿ��� ��ݯ>�P�b�tφ� ��+ϼ��������� Y�k�}�/ߑς�ſ�� �������߱��$�6� H�k�l��ߐ����� ����-�?�Q�2�e�V� ��z�������s����� ��
?���;dv �������%� 9[�<N`r�G ������&/ 8/J/\/n/�/��� ���//?"?4?F? X?/|?�?�?�?�?�/ i?�?OO0OBOTO�Z_ERR m�Z�\OlFPDUSIZW  �0^0��D�>�EWRD ?��U�!�  guest�6��O�O __$_6_�TS�CD_GROUP� 3n�\ �Q��9IFT|^$PA�|^OMP|^ n|^_SH|^ED�_w $C|^COMn@�TTP_AUTH� 1o{K <!�iPendan�BWMn�[�2�q!KAREL:*MoVohmKC}o�o�o�u`VISION SETfP�o�o�v!,rcP>h b������~dCTRL p{M�6��1
F�F�FF9E3��$�FRS:DEFA�ULT[�FA�NUC Web ?Server[�I� �"d�O�D�я������+�jDWR_C�ONFIG q.kU�Bc[�lA�IDL_CPU_kPCz��1B��  BH��MIN���sQ��GNR_I�OuA�B�0�H��NP�T_SIM_DO�ӖݛSTAL_oSCRNӖ �ޚ�TPMODNTOqL�ݛ��RTY��p����` `ENB��sS��OLNK 1r{KxP����ɯ�ۯ������MAS�TEҐy�5���SLAVE s{K�H D��SRAMCACHE/�A�"aO_CFGq������UO�`����CMT�_OPz�ՒJǳY�CLp���t�_AS�G 1t`��A
 �6�H�Z�l�~ϐ� �ϴ���������� �\�	�NUM�CI�
��IPn���RTRY_CNҿ���G_UP_��A����E� ������u)� � 06��م�RC�A_ACC 2v�k[  R��� 1�  j�� 6�� 6���0,�4�4��g 9"�� �2�D���BUF001� 2wk[= {�u��u0����u0pi��u0�n��)��8��I��X���i��x�䉞䘪�䩞丞�ɞ��j�������	���� ���������������Z������������u0�Z�x����!���0��A��P��a���p����������(� ( �V�� ������U$��3��D��S��Ud��s�䄖䓖���u0�l�����Ɩ�Ֆ�s�2��������u{ ��t(�� �����������������t� ������ ����$�) ��)�<�)�L�) �\�)�l�)�|��K *����phȜ������� ��������� ���������������t� � � � �% � - �5 �= �E � M �U �] "e � m �u �s�3��� �.��.�-�@��� .����.����.��� �.���.��.� �#�R%�3�R�$<� K�R�$T�c�R�$l� {�R}��P��P���P ��������� ����������� �����R��#i� #i�+#i�-;#i� =K#i�M[#i�] i��es#i�u���я�2xk[ 46�A��Q�P<�P�D�AՒ���HIS}�zk[� �� 2021-04-21�V ��A�I/_A_ S_e_w_�_�_�_�_�XR��yXCT�_ 
oo.o@oRodovo�o�o���y��;  �L[T�Q18-02-27�_�o�o<�o  T�c,�>Pbt�{LY�3�h5�o��������U�*G�Y�.�sN�2�g1�A��������\��C���BX�Q�``΄hބiC4�D���΄�2��(�:�LM��u�2���q����H<&q��F�:�p΄xބF��A���΄�΄�΄��΄�����rL�� u��`�M�_�q��FՂ Ɛ݂�@��@ђ�`ْ0�@�������Mp� �O_Z: � M�_�q���������˿ ݿ��_;�%�7�I�[�@m�ϑϣϵϣn;�@c�o���%�7�%p5  Z8�c�u� �ߙ߇�������� �)�;�)�M�j�|�j�@|�������ĉ�AdՀ��݀6�d�����X������ -�@L�6Z�O�=�O������ �����Ɛ�ѐ�ⵠ ������͠��ՠ �����	������&� 8�n������݀�� 
���ѐ��� *	�9�L� �&�Z�|����� ��/���/T/f/ x/�/�/�/�/�/�/�d����:/'?9?K?9���#v?�?�?�?�?�� ��?OO*O<ONO`O)�iO�O�O����O �O�OŊ���@݂���@ ��@��~O
�BR�B_ s_�Os��O�_�_���_ ��4Xђ�P���P��
� �P͢�Pբ�P��P	� �P�_oM�_�o�o�o ��$_o$o6oHo�;��I_CFG 2�{: H
C�ycle Tim�e�aBusy>DwIdlzr�t�min={�q�Upvv|qRe�ad�wDow��x�aRqsC�ount|q	Num qr�s�={��`z�!�PROGWr[|:D�0� u���������Ϗ�y%�SDT_ISOL�C  :� ��@~J23_DS�P_ENB  ��>#�INC �}��e�A   �?��=���<#��
�j�:�o u������a��ȟ�+OBK�C,��uU���G_GROUP� 1~�< � �j�Cy.��П?Dxd�m��`Q ������̯������&�Dw��ڙG_I?N_AUTO�Q�>#�POSRE����KANJI_MA�SK��t�KARELMON :(��by���(�:�PL�@~²O��V�X���nŉ���CL_�Ld�NUM0������EYLOGGING��?���U�F��LANGUAGE� :
���DEFAULT� �(LGXq��V��r��d� � 8�pP��`'N6'  ��`ۏ��;��
��(�UT1:\\Ϧ� �ߵ���������� !�8�E�W��(���#LN_DISP �M��x������OCTOL���aD�z@��f��GBOOK �)�=z��qz�z�= �ey�k� }�����������5Ӱs����	-�t�*���/ُ`�+�_BUF�F 2�� 	A�evꂒ �w�����# ,YPb���������/��ZDCS �V�Y�n� ��#Dx^u�/�/�/�/�6$IO 2�B+C cp�/cp@���/ ??*?>?N?`?r?�? �?�?�?�?�?�?OO &O8OJO^OnO�O�O�O~�%ER_ITM��dD��O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogo	�N�BSEV�����FTYP���O�o�o8�ovm��RST��4%�SCRN_FL +2��-@��g/g�y�����T�P�����b�NG�NAM,�`�
�2$U�PS��GIp���U�B�_LOAD��G % �%�ZAD15�O�MAXUALRM��,�� �U�
��H�'_PRM��� !�����C���7���x���P 2�7� �V�	�ol�W� ��{���Ɵ���՟� ��D�/�h�S����� ��¯���ɯۯ�� @�+�d�v�Y������� ������߿��<�N� 1�r�]ϖ�yϋ��Ϸ� �����&�	�J�5�n� Q�cߤߏ��߳����� ��"��F�)�;�|�g� ������������� ��T�?�x�c����������������DBG?DEF ��[!���_LDXDI�SA-��{�#MEM�O_AP'�E ?= �
 $x( �����������FRQ_CFG� ��(A �x'@�E��<[$dA%m$:������*z�/� **:� ����_x&��+/ "/4/a/X/j/�/����/�@�/�/�/�/�',(�/>?�$,?i?P?�? t?�?�?�?�?�?OO OAO(OeOwO^O�O��?ISC 1� �� ����O��)�O���2__V_�O�B_MS�TR ��myUS_CD 1�o�N_ �_J_�_�_o�_4oo 1ojoUo�oyo�o�o�o �o�o�o0T? xc������ ���>�)�N�t�_� ����������ˏ�� �:�%�^�I���m��� ����ܟǟ ��$�� H�3�l�W�i�����Ư ���կ����D�/� h�S���w�����Կj_MK'��]Y�$MLTARM&��-� �3" P�X� METsPUK Ȳ���Y�NDSP_ADC�OLr�& }�CMNmT�� ��FN��|�τ�FSTLI���ǁP ��^'�G��Y?�IԆ�POSC�F����PRPMl��Y�ST��1��[w 4Q#�
�� ϱ�����׿������� 7��+�m�O�a��� �����������E��/��SING_C�HK  ��$M7ODA%��K����DEV 	�N
	MC:��HOSIZEKȰ��TASK %N
�%$123456�789  2}�T�RIG 1��[ l^9n��=YP��5���~�EM_INF �1��`)�AT&FV0E0�+)E0V�1&A3&B1&�D2&S0&C1�S0=)ATZ+fH��:��bA�/�'//K/]/ �/5G Yk�/� ?7/$?6? �Z??~?�?w?�?g/ y/�?�/�/�/2O=?�/ hO�?�OGOQ?�O}O�O �O
__�?@_�?OO )O�_MO�_�O�_�_�O o�_<oNo5oro%_7_ �o[_m__�o�_& ]oJo�;�� ���o��o�o�o�o X�|������e֏������0���NIwTOR�G ?���   	EX�EC1˳s�2y�3�y�4y�5y�C {�7*y�8y�9˳t��r ޔx�ޔ��ޔ��ޔ�� ޔ��ޔ��ޔ��ޔ̒�ޔؒޓ2�2�2���2	�2�2!�2�-�29�2E�2Q�3��3�3���R_�GRP_SV 1ݘ  (7����;=�/";����������?�N?�����
�_Dς��9�ION�_DB���ȱO  �q�y����V�~� Ȱ����ΰ.ΰ/��&�N_   1�������J��-ud1�����υ�PL_NAME !�<��!Def�ault Per�sonality� (from FsD)����RR2��� 1�L6�L�A�<��� d:҉ϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻����������2��.�@�R�d�v�@��������<� ����0�B�T�f�x�����������޲�D����
���P J\n����� ���"4FX '9������ �//0/B/T/f/x/ �/�/k}�/�/�/? ?,?>?P?b?t?�?�?�?�?�?�?�> �H�6 H�b �H\���  �O1M�dC@PO bMFO�O�G@�=�|C��O�M�O�O C  �H__ _2_P_V_t_@�_�f��_�\��E�	`_�_o o�Q:�oA`�@oRodo�vn A�   �i�O�o�Lޱ�o�k�O �o'9$]H�: �R�� 1�4ɴ���R@ � �&�<��p @D��  �q?��s�q?���q�A��6E�z  �q���;��	l�r	 ��@� �0ݰް!� ���p� � �� �F��J���K ��J˷��J� �J�4�JR�<g|v�f0O����@�S�@��;fA6A���A1UA��X{����=�N���f������T;f��X���ڀ��* � ��  �5'��>��p�H���?��?���{#�����ԏur`�f��q{��g�������i�V����(  ����¤��Ȗt柉�	'�� � �I�� �  ���e��:�È(�ß�=���@���߶� <!��� � �  ��qz�˂�r�o�o����ү � '覵��@!�p@�a�@���@��@��C�C�"��"��B�pCz%����@�r��������n���� ���m;a;n�`@����D�u՟ҿ����῀��Q�c�E�Uŕ��w :�W  x�x?�ff�O�Ϙφ*� �P���ˍ�8x�����>��x��q����0�P:�U�7�x0�0���>���|����<2�!<"7��<L��<`N�<D��<��a,h��ߴ��s��s| ҈`?fff?���?&�аT@T����?�`?U��?X�ᒩL� ���t,��t8��wW��� ��ό�w������ �����.��R���!�F�A���=���)����M����HmN� H[���G� F��HZE ~i������ � �oAK���� ����)���/ ��%/7/�j/U/�/y/�/�/��M��"�i���C�/?�/5? =8��`??F??j?��ç�sY��-M�BH"��.��?,�[2�Y0X1�1�@Iܔ=@n��@��@:� @l��?٧�]�? ��%��n�߱����=�=D���0OB@��@��oA�&{C/�� @�UXO�+�J8��
H���>��=3H���_�O F�6��G��E�A�5F�ĮE���O�@��fG���E��+E�?�EX��O�@�>\�G�ZE��M�F�lD�
�p�O�?E_0_i_ T_�_x_�_�_�_�_�_ o�_/ooSo>owobo �o�o�o�o�o�o�o =(:s^�� ������ �9� $�]�H���l������� ۏƏ���#��G�2� W�}�h�����ş��� ԟ���
�C�.�g�R� ��v��������Я	� ��-��Q�<�u�`�r����fB(hA4�̯�h���൘�3��ϩп��!4 ��{����!�0+#8(�:��jbT�f�1E�䴛|�� �ˀ��Ϯ��������JiP��P:�IV c߶�oߙ߄߽ߨف����������9�$��"$<�N��r�����v�H���&��e ,�6�l�Z�|�����n)���������8F
  2 H��6�&H�{�g\Ŵ�&B�!�!� B��0�0A� @�/��$��3���l ^pUgy���$�0� � ��r� T�%
 � �//+/=/O/a/s/ �/�/�/�/�/�/^J�� ��$����4��$MR_CAB�LE 2�$�� � V�TP�
�@{ ?�0F1�?0S��0z Bz C[0�{OM�`B����{�0�#DG��l{??Q6 �� B�� TO
��vr0���5Ų~6q<�|Œ?�8� ��� C� 9h4��r0��2��E�~6�'N�?�?�*�\0�� [@CW@j27��(��{<��2I�/T3�OR˰O �O�O�O�O_�O�O"_ _*_�_�_`_�_�_�_@�_�_oA{+��_ Qocouol�?o�o�o�o�l�*�o** �3OM �%9���z��tc%�% 234567O8901%7u "PRFq{ [@ �{ �{
Lw�nn�ot sent ��jzsW,�T�ESTFECSA�LGRI�gkʝd��t��q
�tG �P�{�"��'�9��K� 9UD1:�\mainten�ances.xm�7��l���DEFAULT~2GRP 2�	z�  p$�  ��%1st m�echanical checkL}6{�6��>�G�H�$r����������{�controller��7��Ic�8�J�\�n����ϑM���{"�8��{ ȡϯH�'�����*�<���C ٟn�����������ҿ����ϒC�g�e�. batt�eryς�W�H	����ϖϨϺ�����Supply g�reasK���{�E�
�<A��g�s�@H�Z�l�~ߐ�� �cabl��߾�g�
7���0�B�T�� ؑ+�����Q����� ������{ $��@�hoo� ������� ����+� O�a�s�) Zl~����� '9 2DV� ��{���� 
//k@/R/�v/� �/�/�/�/�/1/?U/ g/<?�/`?r?�?�?�? �/�??-?OQ?&O8O JO\OnO�?�O�?�?�O O�O�O_"_4_�OX_ �O�O�_�O�_�_�_�_ �_I_om__To�_xo �o�o�o�oo�o3oEo Wo>Pbt��o ��o���(� :���p��_���� ʏ܏� �O�$�6��� Z���~�������Ɵ� �9�K� �o�D�V�h� z���۟������5� 
��.�@�R���v�ů ׯ����п����� g�<ϋ���r����Ϩ� ������-��Q�c�8� ��\�n߀ߒߤ����� �)�;���"�4�F�X� j�ߎ���������� ����m���T���C� �����������3� i�>��bt�� ����/S(�:L^p��	 T~�����/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBOxTOfOxO  ��?�  @� ��O�O�O��O_�_(_�*H_** ���@zO|_�_��_b_�_�_�_�_��!__�_Ko]ooo 1o�o�o�ooo%o�o #5oAk}� �o�oQ���E� 1�C�U����a��� ��ӏ����	��e�w���
�$MR_HI_ST 2��v��� 
 \�$ �23456789C01����P�BR��9���������?� Q�c��,�������t� ��ԯ��ί;��_� q�(���L���˿��� ���%�ܿI� �m�� 6ϣ�Z����ϐ���[��SKCFMAP � �y�*�B�������ONREL  ��v�.�6��EXC/FENB`�
,���y�FNC��r�JO�GOVLIM`�d�v����KEY`�z����_PAN_ظ�����RUN�����SFSPDTY�P��k��SIGN|`�r�T1MOT���o��_CE_G�RP 1�� .�~���O��÷��� a������C�U��y� 0�����f�������	 ��-?&c�� ��t�����Mq(�QZ_EDIT]�(�Q��TCOM_CFG 1�$������� 
�_ARC�_}�`��T_M�N_MODE]����UAP_CP�L/��NOCHE�CK ?$� �� �/�/�/�/ �/�/�/??0?B?T?�f?x?�?�?I�NO_?WAIT_L\�6��NT��$�3z���1_ERR��2�$�6ф�OEOWO�iO�L<юO�O�53 O�C�#M| 1��f?"��A,�:?x��k���µ�B���z��<�� ?����_�O?�7NBPA�RAMB�$���Fg�_yW8ѫ_�[ = ���_�_�S�_ o(oo4o^opoLo�o�o�kxW��o�l}_�n#UM_RSPACE!��b�GQt��$ODRDSP�#_��OFFSET_CAR�_/�v�DIS��sS_A�3 ARK]�OPEN_FILE�p�_���cqPTIO�N_IO�����M_PRG %3z�%$*A�S��sWO��p����Cp쀄����  ;��?֞��g��	 ч�Ȟ����4��dpRG_DSBL'  n�.�J���sRIENTTO�_���C�>�-�A� �rUT_SIM�_D�+ҋBdpV~hpLCT ��=У��O}��d\�_P�EX; ���RAT�;' d�����pUOP �m��pw����� �>�L��$�PAL�2��>`�_?POS_CH�p���`�ZP2��L6߸LA�W����oѯ����� +�=�O�a�s������� ��Ϳ߿���'�9���2��h�zόϞϰ� ��������
��CW�4� F�X�j�|ߎߠ߲��� ������*AAs'�}I5�4�Z�BPG��� �����������&� 8�J�\�n�����a�s� ��������"4F Xj|����� ����0BTf x�������`///_�xW�Y/ k-���c���/�+�/�/ �'>->-�o?�/3?�'tP(7R?H?Z?l?�? �?�?�?&0w��?L�D(4	`<?6OHOZOA:�o<�xO�O�O|�O'0A�  �I !?�O�__�]?>_)_ b_M___�_�_�_u�����O�1���_��� ��$B@ �؄��P� @D�  a?��c�Q?=�a=�D�  Ez0c�:��;�	l&b	 ��@� 0PP_`� �
`� � �� ��b�PH�0#H��G���9G�ģG�	{Gkf���GΈ�K/�o�l�PC�1���`[�D	� D�@ D7g�n�d����  �5��	>(p`�4�(:� B4�Bp{��!=���O	��R��r'a�s0W�Ao�Rҧpߐ��p(  �
�p����_$��U	'� � B��I� �  ���E�F=����f�x���� �<_`� �� � � �ف��8� b__r�WN=��  'N�X(��aOpC�`��`
[pB`Cc5�G� ����@�i����m����G�MuAuN�@@=��*b7e���� 4��X�C����������=�� :�a>�tx?�ff�/į֯h� @��O��8=�3�A�>�� �q"a�J�pn�Px����uancnd؃>�������u<2�!<"�7�<L��<`�N<D��<���,�o��c�� c^��@?fff?��?& �K�@T���2�?�`?U?ȩ?X�B�:� ���'d�Iev�g�� �Zd���ϵ������ ��6�!�Z�l�Wߐߢ� y��߱���aσυ����D���HmN H[���2G� F��M�������� �����(��%�^� _ ���K�����+��� g�*<N�cu������� Β���I={C�Ox�s^?��}����?yç'c�T'sqH�`�xp�ĺ�����:!@I��>}@n�@���@: @l��?٧]/� ��%�n��߱���?=�=D��n/� ���@�oA��&{C/� @��U�/ �+�J8��
H���>��=3H���_�/ F�6��G��E�A�5F�ĮE����/� ��fG���E��+E�?�EX�?� �>\�G�ZE��M�F�lD�
`8?/�?n?�? �?�?�?�?�?O�?O IO4OmOXO�O|O�O�O �O�O�O_�O3__W_ B_{_f_x_�_�_�_�_ �_�_oo-oSo>owo bo�o�o�o�o�o�o�o =(aL�p �������'� �K�6�H���l����� ɏ���؏��#��G� 2�k�V���z��������韤"(�!4��ퟦ����֕3��ϩ� ��!4 ��{:�L��!�0+#8f�x�Z�jb����1E�䴛|� �������"��F�4�J��P޲Px����� ������׿¿��湿����A�,�Q�w�b��"$zό��ϰ����πߴ���@�.�d�R�e j�tߪߘߺ�������)����.��R�@��v��  2 H��6�&H�����\Ŵ�&B##B�  A� @'����@�"�4�F�W���߀�������������$J�� � q�� 9��%
 ��3 EWi{���������* ���b����4��$PARAM_M�ENU ?����  �DEFPUL�SE�+	WAI�TTMOUT��RCV� S�HELL_WRK�.$CUR_ST�YL�OP9T���PTB���C�R_DECSN�i�<,6/H/Z/�/ ~/�/�/�/�/�/�/?�? ?2?[?VSSR�EL_ID  ������j5USE_PROG %eq%W?�?k3CCR��|2��m�7_HOSoT !e!�4O�:T���?-C�?A�/CiO�;_TIM�E�|6�5VGD�EBUGz0ek3G�INP_FLMS�K�O�ITR�O�GP+GA�@ �Lp� [�CH�O�HTYPE
bn�V?P?�_�_ �_�_�_�_�_oo?o :oLo^o�o�o�o�o�o �o�o�o$6_ Zl~���������7��EWOR�D ?	e
 �	RS�@�P�NS��s�JO�!�TEP@}��COL�3���3WLV�0 ���
���5�d�ATRACEC�TL 1����o v�s �����&���DT� Q���S���D � h��t��h� `�r�����	 ��$P ������ğ֟����P�0�B�T�����j���r����������*���j��r��R��  ���ޯ���&��8�J�\�n������R��Ȱk��r�����������Ȱܴ*ܴ	ܴ
ܴ��޿ ���&�8�J�\�n� ��Z�����&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� \������������� "4FXj|�� �����0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_���_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<N` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���_�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/�"/4/F/X)�$PG�TRACELEN�  W!  �_�V �l&�_UP ������!� �!�� l!_CFG M��%�#V!� ���${#�/�(�-�  ��%�"DEFSPD ��,�U!~ �l IN~� TRL ��-��!8�%C1PE_C�ONFI� ��%O��!�$�)�l LID�#��-	~�9LLB 1�~7 ��$B�  B4�3�& �5JOE��/ << T!?�1KPO1OHOjO �O~O�O�O�O�O_�O��O_L_2_T_�_�Z B�_�_�_�_3O�_"o�o'oXo�9GRP �1��<W!@�  �[�V!A�?x�D P�DV�C2�� o�V d,D�i�i�1�0��0Wo)O�1�n#´(s
�kB+pRq�2.hR�V!>'oY>a�����~� =N�=R��3��0� i�T���x����Տ��x����  Dz0�9�V 
 �a��q��� ������ߟʟ��'� �$�]�H���l������)W!
V7.1�0beta1�$�ܠB(�A�?\)A�G��aޡ�>�������ޡA����f�fޢA�p��AaG��Q�Q@�(��`� ��K�]�o����#Apأ�r�0 ����Ϳ߿ڢU!��} ���v�$��H�2ϝ:�KNOW_M  ��%�&�4SV ���9��5 N�����f�9�$�6�Po��"�m�3Mvc����} ��	�"V ���T���PܽԿ���פ�@1ߠ���(�wPV�1MRvcĥ�T~��D��u����OAD?BANFWD�ϡ3{STva1 1ś)��4�5���� �&��� �Q�D�V�h� �������������� 
O.@�dv������2�����V �<%�w`3 !3E��4bt����5�������6//,/>/��7 [/m//�/��8�/�/X�/�/��MA���d�3�'OVLD � ;�ߊ���P�ARNUM  p��?�?��SCHS9 a5
�7�1�9��
EUPD�?�5uTO>�%_CMP_��V0�����'��lDER�_CHKzE��`��ҎFwO�KRSg����pa_MO���H_��O�%_RES_G
���;
8��oi_\_ �_�_�_�_�_�_�_o �_/o"oSoFo9?+U6\F_xo+Ua�o�o �o-S��o�o�o-S  27-SZ Rqv -S� ���-S 0�x��-RV 1���|���@`z$�BTHR_INRg��X1����dc�MASmSp� Z��MNo����MON_QUEUE ������@����$Nq@U�AN8��ۈ�END��_��EXE ��6@B�E���OPTI�O��[��PROG�RAM %Պ%��.��?�TAS�K_IU4g�OCFG �Տ�?ɟ���DATA�����@�@M� 2 �f�(���������@c��΢֯� ����ɣ @6�>�P��b�t�����INFO
���I��䄽�ǿٿ ����!�3�E�W�i� {ύϟϱ���������@��/ߊ������I�� di���@DIT� ���߬���W�ERFLA�V���RGADJ Ή�/A�  ��?�@�w����� ��W�/�?���z��@'<@�9���%?h�0��dm�C�2�%糲+	H�l7�U�2�u?G�A ��t$���*��/�� **:���@������5,�'�����1��1W�9�Q����/�A� o�e�w����������� ��]G=O� s����5�� '�K]�� �/�����y/ #/5/c/Y/k/�/�/�/ �/�/�/Q?�/?;?1? C?�?g?y?�?�?�?)O �?�?O	OO�O?OQO OuO�O_�O�O�O�O �Om__)_W_M___�_ �_�_�_�_�_Eo�_o /o%o7o�o[omo�o�o�oN�	�<��*c Nt����Q�M����PREF ��%�����
��I�ORITY��܆�>��MPDSP������C�U������OD�UCT�������OG��_TG���钍ڂ�HIBI�T_DOA���TO�ENT 1Ӊ�� (!AF_I�NEm� �+�!�tcp+�S�!�udB�{�!iccmj�qXY��ԉ����)� 0��ߟ����ٟ� ��	�F�-�j�Q�c��� ��į��������$B�T�*����%����V����>VӰ
�f��/	���������~��AG�,  ��o�D�V�h�(z��պ��Z뿺�������ϻ�i�EN�HANCE �u�s�A��d�P�7Մ~���������PORT_NUMn�������_C?ARTREP�Ĝ>�SKSTAm��oSLGS��ě��G�T�UnothingX�5�G��Y��{��TEMP �ڑ�e��e�_�a_seiban ���������"�� F�1�j�U���y����� ��������0@ fQ�u���� ���,P;t _������� //:/%/^/I/[/�/�/�/q�VERSI�L����  d?isablej�m�SAVE ۑ��	2670H7K55�(�/E?!@�0G?Y?|�}? 	�8w�$�o�;�?��e�?O"O4OFOTJ�<|?�Ot��5_�� 1�ě20�@r�e�O�O��g�pURGE�B掘�WFP�p�����W�3T�ѯ�W�RUP_DELA�Y ���&UR_?HOT %!vz��?߳_DUR_NORMAL�X���_�_�WSEMI�_�_;o�q_QSKIP�C�|��Cx�/�o�/�o�o�o �m}�o's�o!3E iW���w� ����/��S�A� c�������s�я���� ��ߏ�O�=�s��� ��]�����˟���>SRBTIF4T��RCVTMOU������/�DCR��C�^i ���aB.&�B����B'�w@�q�y@�)ݹ�4�m�,���e��p]2�)�é�9��oݯ�o<2��!<"7�<L���<`N<D��<��ɫ0�ׯ@�Q�@�u������� ��Ͽ����)�;��o�RDIO_TYPE  �M1�G��ED�T_CFGg ��KbBHS�E��Xa2�� �ȸ�����.�  �үD�/�h�S��ϙ� (o���o��ӟ����� ;�)�_�M��m�ߴ� 9�{��������%�� 5�7�I��������� a�������!E3 i�����a�]� ��A/e� ��mG���/ �+//O/qv/�/G/ �/C/�/�/�/�/�/'? ?K?m/r?�/S?�?�? �?�?�?�?O�?!OW?�}?nO;���INT �2�Y���_�G;� �O�K�+��OX�f�0 _[3O6_ 'OF_H_Z_�_~_�_�_ �_�_�_o�_2oo*o hoVo�ozo�o�o�o�o �o
�o.@&dR �v������ ��<�"�`�N���!��EFPOS1 1��d�  x \O҉���O����+� ŏ׏�r�]���1��� U�ޟy�۟���8�ӟ \�������-�?�y�گ ů����"���F��C� |����;�Ŀ_���� �����B�-�f�ϊ� %Ϯ�Iϫ����ߣ� ,���P�b����Iߪ� ����i��ߍ���� L���p���/���� e�w�����6���Z� ��~��{���O���s� ���� 2����z e�9�]��� �@�d��� 5G���/�*/ �N/�K/�//�/C/ �/g/�/?�/�/�/J? 5?n?	?�?-?�?Q?�? �?�?O�?4O�?XOjO OOQO�O�O�OqO�O �O_�O_T_�Ox__ �_7_�_�_m__�_o o>o�_bo�_�o!o�ox�oUc��2 1崏 ^opo�o(LRop �/��e�� ��6����/��� {���O�؏s������� 2�͏V��z����9� K�]���������@� ۟d���a���5���Y� �}������ů��`� K������C�̿g�ɿ ϝ�&���J��n�	� �-�g��ϳ��χ�� ��4���1�j�ߎ�)� ��M���q߃ߕ���0� �T���x���7�� ��m�������>��� ����7�������W��� {���:��^�� ��ASe�  �$�H�li �=�a��/� ��/h/S/�/'/�/ K/�/o/�/
?�/.?�/ R?�/v??#?5?o?�? �?�?�?O�?<O�?9O rOO�O1O�OUO�O�o�d3 1��o�O�O �OU_@_y_O�_8_�_ \_�_�_�_o�_?o�_ co�_o"o\o�o�o�o |o�o)�o&_�o ��B�fx� �%��I��m���� ,���Ǐb�돆���� 3�Ώ���,���x��� L�՟p�������/�ʟ S��w����6�H�Z� ��������=�دa� ��^���2���V�߿z� Ϟ���¿��]�Hρ� ϥ�@���d����Ϛ� #߾�G���k���*� d��߰��߄���1� ��.�g���&��J� ��n�����-��Q� ��u����4�����j� ������;������ 4���T�x ��7�[� �>Pb���!/ �E/�i//f/�/:/��/^/�/�/?�OT4 1�_�/�/?�? m?�?�/�?e?�?�?�? $O�?HO�?lOO�O+O =OOO�O�O�O_�O2_ �OV_�OS_�_'_�_K_ �_o_�_�_�_�_�_Ro =ovoo�o5o�oYo�o �o�o�o<�o`�o Y���y� �&��#�\����� ��?�ȏc�u�����"� �F��j����)��� ğ_�蟃����0�˟ ݟ�)���u���I�ү m������,�ǯP�� t����3�E�W���� ݿϱ�:�տ^���[� ��/ϸ�S���w� ߛ� �Ͽ���Z�E�~�ߢ� =���a����ߗ� �� D���h���'�a��� �����
���.���+� d����#���G���k� }�����*N��r �1��g����8?045 1�;?��1��� ���/�/Q/� u//�/4/�/X/j/|/ �/??;?�/_?�/�? ?�?�?T?�?x?O�? %O�?�?�?OOjO�O >O�ObO�O�O�O!_�O E_�Oi__�_(_:_L_ �_�_�_o�_/o�_So �_Po�o$o�oHo�olo �o�o�o�o�oO:s �2�V��� ��9��]��
�� V�����ۏv�����#� �� �Y��}����<� ş`�r������
�C� ޟg����&�����\� 寀�	���-�ȯگ� &���r���F�Ͽj�� ���)�ĿM��q�� ��0�B�Tώ������ ��7���[���Xߑ�,� ��P���t��ߘߪ߼� ��W�B�{���:��� ^���������A���xe�K]6 1�h �$�^����� �$ ��H��E~�= �a�����D /h�'�K� ��
/�./�R/� �/K/�/�/�/k/�/ �/?�/?N?�/r?? �?1?�?U?g?y?�?O �?8O�?\O�?�OO}O �OQO�OuO�O�O"_�O �O�O_|_g_�_;_�_ __�_�_�_o�_Bo�_ foo�o%o7oIo�o�o �o�o,�oP�oM �!�E�i�� ���L�7�p���� /���S������� 6�яZ�����S��� ��؟s����� ���� V��z����9�¯]� o�������@�ۯd� ����#�����Y��}� ϡ�*�ſ׿�#τ� oϨ�C���g��ϋ��� &���J���n�	ߒ�x���7 1��?�Q� ��	���-�3�Q���u� �r��F���j���� ��������q�\��� 0���T���x����� 7��[��,> x����!�E �B{�:�^ �����A/,/e/  /�/$/�/H/�/�/~/ ?�/+?�/O?�/�/? H?�?�?�?h?�?�?O �?OKO�?oO
O�O.O �OROdOvO�O_�O5_ �OY_�O}__z_�_N_ �_r_�_�_o�_�_�_ oyodo�o8o�o\o�o �o�o�o?�oc�o �"4F���� �)��M��J���� ��B�ˏf������ �I�4�m����,��� P���럆����3�Ο W����P�����կ p���������S�w����6����߷�8 1���l�~���6� !�Z�`�~�Ϣ�=ϟ� ��s��ϗ� ߻�D��� ���=ߞ߉���]��� ��
���@���d��� ��#��G�Y�k��� ��*���N���r��o� ��C���g������� ����nY�-� Q�u��4� X�|);u� ���/�B/�?/ x//�/7/�/[/�// �/�/�/>?)?b?�/�? !?�?E?�?�?{?O�? (O�?LO�?�?OEO�O �O�OeO�O�O_�O_ H_�Ol__�_+_�_O_ a_s_�_o�_2o�_Vo �_zoowo�oKo�ooo �o�o�o�o�ov a�5�Y�}� ��<��`����� 1�C�}�ޏɏ���&� ��J��G������?��ȟc��ҿ�MAS�K 1����0�>��XNO  ��=�C�MOTE�  _�  ��_?CFG 휭���PL_RAN�G������٦OW_ER ������SM_DRYP�RG %��%���I��TART ��	�W�UME_�PRO&�8����_�EXEC_ENB�  ����GScPD��ΰָ�gTDB��RM���I_AIRPUR� ��m�p��MT_�T������OBOT_ISO�LC]��l�̥ȥ���NAME ����OB_O�RD_NUM ?�	�i�H?755  ��@��R�d��PC_TI�MEOUT� x��S232��1��`�� LT�EACH PEN�DAN�б�С��������Ma�intenanc�e Cons�������"�ߒ�No Use�����@��R�d�v�����NPqOf���С�����CH_L������	���!�UD1:1���R�VAIL!ц��������SPACE�1 2�`�
��ХЩ�巓ΦТ��m���< ���?�Y�Y��� KlC�|������ ���%<�Q rY`�d����� �Y)/@/�U/ v/]/�/����� �//7/-?�/Q?r?�? k?�/�/�/�/�/�?? 3?)OJO	O_O�OgO�O �?�?�?�?�?OOAO 7__[_|_�_e_�O�O �O�O�O�__=_3oTo ou_�oqo�o�_�_�_ �_�oo)o/Moe �]o�o�o�o�o �%G=�^���� {���������!� S�9����o���g���t���2��� �� ݏ����%�W�Z���@:�������Ưǟ3ڟ ����"�ԯF�x�{����[���ҿ����4 ����1�C���g��� ���|��������	�5�.�@�R�d�߈� �Ͻ�ߝ������)�*�6=�O�a�s߅�7� ������$���5��J�K�7^�p���� X�������E���5V-kl�8������� ��y�� f V�wN��G �N� �ń
�7 �  �/ /1/C/U/g/y/����-���/m�/ȁd 0�/2?D?V?h?z? �?�?�/�/�.�:�?�; O??�?ZOlO~O�O �O�O�?�?�?�?O_ 5_(O:O�Oz_�_�_�_ �_�_�O�O�O _"_4ow `� @Ȁ�me�/{oW__Y�a�U Do�o�o�_�j�o�o1 CaI��gq �������Q� c���7�i��������� ��Տ�ُ�\
�ol���A��*SYS�TEM*�V9.�10185 ��1�2/11/201?9 A �� ���r�ӓSR_T   � $Đ�ENB_TYP �  $RU�NNER_AXS�� $HAND__LNGTH�`��THICK��FL�IPґ�`$IN�TFERENCE|��IF_CH���I֑$�9�IN�DXD�ĐG1POS   W�\N�`�ANG`�x�w_JF��PRM`�� 	�RV_D�ATAƑ  �$��ETIME�  ��$VALU�����GRP_ �  ��A�  2 �S�Cő	� ��$ITP_�� �$NUMڠOU�ِ	�TOT�
�D�SP!�JOGLI�M� $FINE�_PCNT@�CO|��$MAX��TASK@�KEP�T_MIR=�]�P�REMTq�}�AP9LD���_EX���`���t�@��PG��BRKHOLD�t!��I_�  ڲ�@���P_MADyE�w�BSOC��MOTN�DUM�MY163�SV�_CODE_OP�M�SFSPD_O�VRD��R�LDlL�O�ORZ�TPӐ�LE[�F!�[�:�OV=�SF��ᐓ�T��F��A�a�UFRA���TOOL@�LC�HDLYW�RECcOVK��:�WSs�:��=�ROM��I��_�ڐ @��S���NVERT�O�FS;�CǠD�FW�Dt���p��ENAYB��7�TR��`����E_FDO��MOB_CM���B-�BL_Mi�]��Ҫѽ2S�VSTAA�G$UP�����G����AM����а��%�f �_M��A�AM�<A�1�T$CA0�,�uD�7�HBK����L�IO?�[�I>Q�$PPAO�{��`��s��s�1�DVC_DB��F���� 쑼��A���1��%����3��+�ATIO"� �h�K�U��/�,/�P�ABF�T֒E��G�Ԛ���E�:�_A�UX�SUBCPyU�G�SIN_7Ј����P�1������F�LA��ݑHW_C�1���j�����$�ATR���$UN�IT�����AT�TRI���G�CY{CLC�NECA!����FLTR_2_�FIR�TARTU�P_CN`Ӷ�SIGNO�LPS�2�1�o_SCTz�F_��cF_��t��FSF����CHA��[�8��O��RSD/���/�P��s�_T��P�RO�|�p�EMP��=��T���ܐx���'DIAG�?RAILAC��p�M�LO��'�4&�PS-�@� i�+��%�PR��SB� � �C�� �	$�FUNC��~�RINS_TB�0��=�o�RA���`�7��a�E��W�ARq�8�BLCU	R�$A+	((�DA��G(#%L�D=�?�h�o#��to#TI��%�ܐ�$CE_RIA�_SWA�AF��Pb^��#��%T2\sCK��CMOI��>�DF_LE�_��PD�"LM��FA>�HRDYO��E�RGt H� z���O >5MULSE� ����0��$JW�J�rǂ�FAN_A�LMLV�Î1WR=N�5HARDאO�_O,� �2�1S�TO�Ƶ_���A�U��R�(���_SBR���5.�J���|�CMPINFڐ���-De!8CREG�@�NV0l�$�۱DoAL_N��FL����$M 2��7%�ܐ�8�ECM-�N0�Y����G����SP$R�$Y���Z����ۡ��o� ���EG!`
�?�
QAR�0�'��20�U3 ��AXE�$�ROB!�RED&!�WR�߱_i]�CSYܰDQᰋVS�W�WRI�V��ST�R �)��f�E�� Ġ&To�1�B�P1�r�V5c�OTOHA9Ġ�ARY�b0]�ΡR�FI��h�?$LINK�!��~3a$EXT_�S�1�%U6�[aXY�Z�2ej7sfOFF�9�2bZbNh`B���d�����cFI �g�A�7Ĩ9�_JL�¢d�?c�h��0�T�[8�US"��B	qL2ArC7 ���DUO�$V9pTU�R�0X�#zu!a(BX�P,�)wFL[`��@�0P�p|e�Y30�Gѯ 1ĠKF�M�'�3��s�����a�ORQ.���x ��s��m�� �H��8,�_A]�OVEd���Mh l��C~��C~��B }��0{�B�|���{�~� �h� ��e�u����� l�v�e�����C����.�ERK��	tE�Ъ��E�A�ܐ��e� gN!K�N!AX�¢N!���4b�� 0��Z1��o��`�� r`���`��:p��qp��1�p��:0��:0��:0 Ǚ:0י:0�:0��:0��:0�:0'�D�8�D7EBU��$��30(�N�VbABNL��t�^�VA�� 
 ����+���7�0�7� o7�a7�ra7��a7� :q7�qq�$Fp�"ۂ�cLAB�b)�����GGRO: )r�<*�B_,��Tm��`�0���*���1�AND�pt�:�+�_e=��1Y� *��A�Pm�!|Ȍ- ^`NT�0ӟ�V�ELل��L����SERVE���@� $�`�A]!��PO@ҹ ��`����ÿ!�@  �$�TRQ�r
� �tR
���"2��q I_ 	 ql���[ERR�b�oI,��لr�TO	QلրLHP���R��� G��%Ha��  � �REP  
 �,��#�=�݁RA~�� 2	 d���s��@��� �@$r�� ���@��OC?!� � d�COUNT��Q ��@FZN�_CFG	� 4��aF3T������ܣ�q ���xR��C �(�M��g2��0Ճ{����FA� ��&��XdP�����$SQ��G�dQPB��@�HEL}@Y�� 5pB_BA�S��RSR`F�"^SS��!M�1��M�U2p�3p�4p�5p��6p�7p�8��@�R�OO�p��V ]`NL��ALsAB��FN�A[CK�IN�Tg CU�0E0� 	_P�Udq�2ZOU��P��aH-�֨ �P��T�PFWD_KAR�w�iAf�RE��$0P8/`U!w�QUE`I  e�Up�r�0�1I�0��-�[`S��SF[aSE�M3��A�0A��S�TYSO� 	�D�I�}����!_�TMuCMANRQ�L[`END�t$�KEYSWITCaH^s.�HEUp�BEATM�PE�PLEv�����U�rF�sS3DO/_HOM� O�1 EFA�PR�a�vQ�P�EC�O01c��яOV_Mr� � IGOCMGt�A�	Pv,�HK�A DXa$bG��U^ҹMP��W�WsFORCfCW�AR 2P�.�OM>P  @��c*�0U�SP3P1�&�@��$3�&4�C"�Oʃ L�"��aHUN�LO9 \�4ED��1  �SNP�X_ASZ� 0Ί@ADD��$�SIZfA$VA����MULTIP���.3� A�! � $H	/0�$�`BRS}�ϱCrТ6OFRIFu��S� ص)��0NFOODBU�P~��5�3�9���AfIA�!$V�y�x��R�SN��@ �3 L0��TE�s8�.:sSGLZATAb�p�&o�sC᳍P[@ST�MT�q�CPP�VByWe�\DSHOW�Env�BAN�@TP�`��wqs8��s8��r"�V�7�_G�� :p$�PCD �7���FBZ�!PXSP� A �U��VDP���� �W�A00 ^�ZR� bW� bW� bWT� bW5`Y6`Y7`YU8`Y9`YA`YB`Y@� bW��cV�@bWF`X 7�$hlY(@$h�Y@@$h��Y1�Y1�Y1�Y1��Y1�Y1�Y1�Y1�i1i1"i2_Y2�lY2yY2�Y2�Y2��Y2�Y2�Y2�Y2��Y2�Y2�Y2�Y2*i2i2"i3_Y�pT�xyY3�Y3�Y3�YU3�Y3�Y3�Y3�YU3�Y3�Y3�Y3iU3i3"i4_Y4lYU4yY4�Y4�Y4�YU4�Y4�Y4�Y4�YU4�Y4�Y4�Y4iU4i4"i5_Y5lYU5yY5�Y5�Y5�YU5�Y5�Y5�Y5�YU5�Y5�Y5�Y5iU5i5"i6_Y6lYU6yY6�Y6�Y6�YU6�Y6�Y6�Y6�YU6�Y6�Y6�Y6iU6i6"i7_Y7lYU7yY7�Y7�Y7�YU7�Y7�Y7�Y7�YU7�Y7�Y7�Y7iu7i7"d �@�P�U� ��߰e�
FQ�2��/ x #�R�@+  ��M��R9� ��Q_+�R����(є~ ��S/�C�D��^�_U�0i��"YS�L���� �  L5Bj��4A7�D��<��&RVALUj�% �x1���F��ID_YL�3��HI��I�"?$FILE_L!��i$�n0��SA�� h	�M�E_BLCK�Z�uA>c�D_CPUs�M0@s�A0u�$�6�E@YZ@�FR  � �PW-����0��LA�AS�������RUN_FLG�� �� ���v�!���!���HF ��C����AT�2x_LI�" w ��G_O�}� P_EDI�"c [���c�k��9��nє0�!�TB{C2LT �Q@` �(0�!c�FT�\��	TDC�A4�z���M�������T�H�0�!�#�$�Rx��0e ERVE�F�	F�5A�� ��  X -$q�LEN�~�	q��) RA� 2��W_�?���1q��2��MIOk�5S�0 I. �Z�����q���DE<�1LACE,":��CC3Z¶_MA�20>>TCVEfTXg
�|
@8R1Q�1QJ%A-UM���J>JPR�}�2�`�@0P	0JKVK�A.)A.5A#�J�AF2JJ:JJBAAL2h:�hbAAf5#� NA1��XB G�L��a_�A�0����CF62�! `	�GROUP��vA�2$QN��C�3~�REQUIR1��0EBU�3m��$T 2 *!n�&8��50��" \� ��oAPPR  CLG��
$t�Ng(CLOD��w)S��)
��.u6# ���M �C 8� 2�$_MGA� �CLPN��(� R �'B{RK�)NOLD�&�@RTMOb�:
=�%Jb�4Pj  :�  B  �  �  6W57W5hA�m��$� "���A��7)A�3PATH �7�1�3�1���3� / 9#\�PSCA�� 7lh"�!INp�UC����0@C:PUM9HY���� @A��L�[J��0[Jq0[@PAYL�OA7J2L�R'_AN��CL�ЦI�A�I�A�%R_F2�LSHR@��ALO��D~A�G=C�G=CACRL_��-E P)G�Dr�H��G�$H�"^NRFLEXj#��J��% PT"�����E�W��jQp�& :}��� �W�T���� ������F1 �QEeYg������(�bE2DVhz ����`x}t�� m`�x���Q	T�w^qXF���d �h%.�x1CUg ktb�����vY�BJ�' ���`��	/���ATrf!� EL�`(�D�#(�J/ &* JE0C3TR)AmaTN��@��'HAND_VB�G�jQ���4( $��pF2�&���S�W�!	��&)?� $$M�@�) !��!�1�#p��E2�A���@�&��<��-QA�,���*A;A;PG��+���*D;D;eP�0G��ݩST�'h�9�N8DY� e �&(�O��@r��G�Q �G�A�G�t`�5P_5h5q5z5�5�5�5t�2�J��* ��T�2 �a㵙!�OASYMEZ� BF)K� L�A$O_B� X5@HD2=4ĸ�ROdOvO�O�CJ�LR0�J�ø���Id_VI��xؙ#!�V_UN���6�W��AJN�|� N��LR�U_ԃ�]� @$YR03_E_���[T�cS�"��HR���a+���}P]"DI0�#O#�2��,) g�V�I9�AV1S P�s`^�^�v`���`� - � ɑME�a��y���`�T�PT��Հ�0����V ��������T��� $D�UMMY1q1$�PS_p`RF2` � �0���PFLA��YP���$GLB_T��1����]!�P�`q�}�. �XT '�1ST��* SBR�0M21�_V&"T$SV_�ER�@O��w��C)LK�w�A�`OS� ��GL�EW�/ �4���$Y��ZB��W���AœAz�9B ��U��0� �pN���$�GI��}$�� �/�0�����1� L���}$Fz��ENEAR�`�NwcFd	�`TAN9Cwb�1JOG&`H0� 2t�$JO'INT�"� iP���MSET�3  "EJ�a�S����1��4� �n`U�a?�* LOCK_FO�@Б�oBGLVt�GLTEST_XMj N�EMP� &"2I�� $U�P��9`#20* ��X1#̐4� X/y�CE�&�y $KAR$qM>%�TPDRA����VEC`�� I�UX2]HE T�OOL9c�V8dR�E�IS3�U�6�z1m`ACH� / 3��O@����3g��% SIZ"  @�$RAIL_BO�XE���ROB�O)?���HOW�WARVQH!��!ROLM�n%ԁ$"p�6 a`�0O_F��!��HTML5��)AͲ��!�15���R�O�R6��"1`�� �ӽ�O�U�7 d��T/�`�J�$�� $PIP*N�p�6"!`�X� �PCORDEaD� 
@� a XT*0�) � �O`� �8 D 0�OB |�N�� �7v1��/�v2܊�P�SYSv1ADqRO� ��TCH�� 9 ,�pENT	�QA_�4�݁@�u�PVWVA~|�: � �����PREV_R�T��$EDIT�(FVSHWR�Pc�G@�b���D���O�^DW�$HECAD����x@��0C�KE����CPSP]D�FJMP�0L�2iPR�`;�;~0{Q��6I3SO�C��N�E�P���TICK�9c��M�Q��CH=NY�< @�0�AᅗA_GP&V-&�PgSTY�2!LOK��Ȑ�D"R�P= tk 
#@G�5%$A�=c�SE�!$@D�9`���M��P&�&VSQU�,e�яTERC�ਁ6�S�>  o�� �p��q�``O����F{`IZ����PR\0�Db�A0P9U;�Te_DOi�0�XS� K�AXI4s`�#]UR��c@P�O P�6���_��2ET�bP�0	�%rPF	�sPA����9'[) �z�PR��?l�P �!���/u�Ay�/u *�/s8�/sH�uuj�uu z�uu���u�}���u�|$���yC
��}C�}��p�ϧϹ��SSC3�� @ h��DS�4P���SPJࡅA	Tx� �UaP�B��ADDRES�B�3@SHIF�O_W2CHO��1IR���TUR�I�� �A�"CUSTO��d x�TV�I�>�B�2��8c�
�2
rV1da~�C \a�8�rPC�a�P��C��b�bR�6����TXSCR�EEx2D��QT�INA��# Ӕpq�a��ٰE T�A ��8b�1��n� ��a�28�b�/@RROS�~ `�0�@�o� UE�DGF ���1
�S��N�1RSMPwgUe00�P抡�S_��@=Ú���ȧ=õaC����� 2E��U�EմGD���D`G+MT��Lp��a~��O�
�BBL_r W��~�H �rPjJ�O��V�LE��a�N �`�RIGH�j�BRD��ہCKGR����Tf0����WIDTH#T@�b�)!��)�UI&� EY��}�I
2� �m VR6 @aBAC�KTQ�Ũ���F�OS1�LAB_q?�(��I �$UART!E���ް��H@�� J 8��~ _wA�h�R���s�(��u�U�O�~�K�P����Uv���Ry!LUM�ØfՀ'ERV!1R�Ph �5L���`GEI�O��`l2�@LP��bE�Pf�)%�v�3؆�3�T  2�50�60�70�8��R��?`h ����j !�S�PKݱ�USR��M <�a���U(�FO\�PRI�am  ����TRIP2!�m�UNDO;�N� �P �ye`!xe�q�O�`�P Oc�\��CaG PT� �T��^�OS��s�R �`F�J��Z�P���� ����6Th�PU�Z�Q���ã�5UJ�OSFF([�R_���=O)� 1P���Z;�Q��GU�1P:���"V�Q�`��SUB86R���SRT��taSR}� #cOR N��RAU(p��T����7��_&@�DT |�1p�8OWNM��4�$SRCQ�Ҡ�PDx(&rMPFIMT|��`ESPPab� ���eA�������A@n
�U `��WO[pr�4a�PCOP��$�`O�_- b�,1�WA3@CF� � Z���@l"+�� V�SHAD�OW�`��_UN�SCA��ʴD�GD!�1EGAC<�8�x�VCWp`>
�W� ,"w16�S$NER�cȷQ#+�C0cDRkIV6f�a_V/P��@m D��MY_UBY��kyV��UR��P�eA�h "�P_MT"LZkB�M]�$�@DEY��3EX7�^��MUb�@X]�V$��US���`�_R��R��
��R��QG�pPACIN�A�PRG�$�"��"��"ң�RE}�遚�:�H�"@�X �� G�P���� �IR��@Y ��?�ӱ��	�qa�REb#SW� _A$�!<�W#B`O��ہQA�^3/rE��UeP��;�6HKjRZ��v:�P&q[0%��3EAP�7� j�^5۰�IMRCV
�[ U��OvPMj�C���	�2��#�2REF 6�F�6�1M0���c50 ���:FAJFAKhE�6��?_ �:�H�;�pS ��N'�aaQ�I�\ �GR�ӵ`����POU4W�"V�k W 5U�2���$Ԑ��C`,�Y`��U�2Q{�ՀULj��Z_ CO~��[H EPNTZ�Th@�U���V�ђSQPL���U#�U���W����VIA_���] ̈́�`HD����$�JO��6��$�Z_UPL�W�Z�|pW!e�QPSp�0�_{LI��$EPEQ ��k�a�QǑ΁��΀��@\m�^� 0贃�a� ��CACHLO:A�d�aI оi��� 1CI`MI�FHa�eT�p�f�K�$HOj��`C'OMM���Ot�w�WӲ�S&�T7 V�P�"@�mr_SIZwtZ� rx!asw�v��MP�zFAI!`5G�4�`AD�y��MRET�r|wGP���> & �ASYN�BUF�VRTD��%�|q��OL�Di_��A�W��PC���TU7#�`Q{0	�EwCCU�(VEM� x�e���gVIRC�q�9�!���%�_DEL�A�#&Q���AG:5�RK!XYZ̠��K!W1��8A��򱦀TN8"IM߁8���|���eGRABB��Yb"��e�_����LAS��<��a_GE�e`u�&��;���T/S&N` ���%aI���"ņ�BGf�V5��PK� ǆ�aWGI��N#�`2�񐂑�`�qq�a+�aS��p�fN:��VLEX��b�����;��Nq��I? �-|�� |�.$�3k��- 
�"c��b�t�Ŀ�\�a�ORD����p��w�RN�d $MPTIT� �C���F�VSF����e�  -�[�QK UR���VSM!�f+���ADJ�N%�P;ZD>�g DƨBa�AL+`�p�AbPE�RIs`��MSG_Q9�$}q�u���b��h+�"�g�J`�^3p�XVR#�in��b�T_OVRi��_�ZABC��j�"(;�s/@
1Z]�#�k+�=$L�-B��1ZMPCF��l�H���A����LN�Kc�
����m $,q�0�įCMCM� C�C����p4P_A+A'$J����Dbq� ��h �h ����
D��F�UX���UXE]!f��	�]��]��oс�oё���FTFpsQӾ�r1 �Zb�n {�}�����uYJ`D�� oY��R�pU�$HEgIGH�#"�?(MP��.A�P���Dp g� EX�$BQPxx �SHIF�s��RVI`F��/B|�0�C`�dTF {"��������WuD��T/RACE��V�A��� PHER� �q ,MP�)�;�m��$R�!p�� ����F�' S�6�S��F��  S�x�2p������s���r�D����	��U�C��ADC���l6�R  d�� Z@D �Qx0C����l�Xl0�| �6�9V��@ 2F���_� D� P�� ���	�	F�,:$ ZH~l���� ��� //D/2/h/ V/x/�/�/�/�/�/�/ 
?�/??.?d?R?�? v?�?�?�?�?�?O�? *OONO<OrO`O�O�O �O�O�O�O�O__8_ &_H_n_\_�_�_�_�_ �_�_�_�_�_4o"oXo Fo|ojo�o�o�o�o�o��oF��$SAF_DO_PULSC� G��k�$qp���|�k���5qR ���`�X{P�S�%S�
������s��tq ��� �����*�<�N��`�r������ � ��2��tqtqd��������rs�� @������*�܉��� � 6��_ @J�TY J����������T D��������)�;� M�_�q���������˯�ݯ��~�����M�_�$��sR�;��f���p����
�t���Di��q��  � ����R�q|u lq���%�7�I�[� m�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w������S��G������ �0�B�T�f�x�� ������������" 4FK��b0E�ҳ D�ܽ������ '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?��?�?�?�? �?�?�?	OO-O��QO cOuO�O�O�O�O�O�O Lz��!_3_E_W_ i_{_�_�_�_�_�_�_ �Yoo,o>oPoboto �o�o�o�o�o�o�o (:L^p��@�����ø�� Ǔ�6�H�Z�l�~��� ����Ə؏���� �2�D�V�d�#�m���.�������i��	123456�78ݲh!BO!ܺTz1!���
��.�@�R�d� v�������"�ïկ� ����/�A�S�e�w� ��������ѿ����� �)�;�M�_�qσϕ� �Ϲ���������%� 7����m�ߑߣߵ� ���������!�3�E� W�i�{��L߱����� ������/�A�S�e� w��������������� +=Oas� ������ '9��]o��� �����/#/5/ G/Y/k/}/�/N�/�/ �/�/�/??1?C?U? g?y?�?�?�?�?�?�? �/	OO-O?OQOcOuO �O�O�O�O�O�O�O__)_;_BS��]_o_��?�_�_�_ԚC�z  Bp�z  � ��2�� �} �X
g�/  	��R2U_<o�No`oro�l��\� +o�o�o�o�o"4 FXj|���� ������oB�T� f�x���������ҏ� ����,�>�P�b�t����������Qa�R�<Ք ˕a  ��������#a#at  ��P#�;���`�$S�CR_GRP 1��*P�3� �� ��R� �U	 /������� ���Qԑ�U������ٯ8ǯ ��]�`��C�,����m��C�����lLR M�ate 200i�D 567890�!`LRM|� 	?LR2D ���?
1234��ЦA�d��hbճ����}�ݣ}��cԑ����ѡ�	j4�F�X��j�|τ���H���Ē�}���į@������̦<��1��@A���e��WV��Vh`�,R��  -���B��Pư߮���Ԫ�A�P��  @��0�ժ�@����� ?4���H�P'������F@ F�` Q�Y�P�}�h���� ���������ʩ������J�5�G�Y�k�B� y������������ =(aL�p���o�
'�����W�`�.4�@4�>'�1U4̧@��n�PȄ����ݣT_��A���ߒ���aĲ�1  
/1/C/Q*!f(r/$�/S/�P�#
b�/ �/�/� ?�/$?,4]��ECLVL  ��1����>1L�_DEFAULT�F4������0Z3HOTST�Rf=�z2MIPO/WERFE0�Ur5��4WFDOg6� r5=2RVENT� 1M1M1�3 �L!DUM_E�IP,?H�j!?AF_INEf0+O�3D!FTOZN�!O~O!�ϣO ��mO�O!RPC_OMAIN�O�H��O�_�CVIS�O�I��_b_!TPUPP�UY_IdQ_�_!
�PMON_PROXY�_Fe�_�_uR��_Mf�_Fo!R?DM_SRVGoI9g5o�o!R���o�Hh�o�o!
�@M�oLi�o*!R�LSYNC+Qy�8v!ROS� O�|�4e�!
�CEwPMTCOMd�Fk��!	�rOCONS�Gl��Z�!�rWASR�CaoFmI���!N�rUSB��Hn�� �O�Uc���?�d��+���O���s�П87R�VICE_KL �?%�; (%SVCPRG1ןD�	�2�$��3G�DL��4o�t��5��D���6��į�7� ����/�*�97�<���od������ 9����a�ܿ���� ���,��ٯT��� |��)����Q���6� z���6����6�ʿD� 6��l�6�ϔ�6�B� ��6�j���6����6� ��4�6���\�^�
�ܟ ���������.��� ���8�#�\�G���k� ��������������" F1X|g�� ����	B -fQ�u��� ��/�,//P/;/ t/�/q/�/�/�/�/�/ �/??(?L?7?p?�_DEV �9�UT1:|?~�0GRP 2
�5��0�bx 	_� 
 ,�0x? �?�2�?OO@O'O9O vO]O�O�O�O�O�O�O �O_*__N_5_r_�_ �?�___�_�_�_o�_ &o8oo\oCo�ogoyo �o�o�o�o�o�o4 �_)j!�u�� ������B�)� f�x�_����������� ��M�,��P�7�t� [�m�����Ο���� �(��L�^�E���i� �����ܯ�� ���� 6��Z�l�S���w��� �����ѿ���2�D� +�hϿ�]Ϟ�U��ϩ� ��������@�R�9� v�]ߚ߬ߓ��߷��� ����*��N�`�G�� k����������� &�8��\�C�����y� ��������C���4 F-jQ���� ����B) fx_������ ��/,//P/7/t/ �/m/�/�/�/�/�/?��/(??!?^?e3d �e6	L?�?�?�?�?0�?�?OK%�O5O<C���NA�1NE ^OlGVO�OzO�O�O�O �I"O_JI�O4_"_X_ F_h_j_|_�_�O�__ �_o�_0ooToBodo �_�_�o�_�o�o�o �o,P�ow�o@ �<�����(� jO�����p����� ��܏ʏ �B�'�f��� Z�H�~�l�������؟ ���>�ȟ2� �V�D� z�h�����ůׯ���� ����.��R�@�v��� ��ܯf�п������ *��Nϐ�uϴ�>Ϩ� ���Ϻ�������&�h� Mߌ�߀�nߤߒ��� ����.�T�%�d���X� F�|�j�������� *�����.�T�B�x� f�������������� *P>t��� ��d���� &L�s�<�� ����/T9/K/ /$/�l/�/�/�/�/ �/,/?P/�/D?2?T? V?h?�?�?�??�?(? �?O
O@O.OPOROdO �O�?�O O�O�O�O_ _<_*_L_�O�O�_�O r_�_�_�_�_oo8o z__o�_(o�o$o�o�o �o�o�oRo7vo  jX�|���� *�N�B�0�f�T� ��x�������&��� ��>�,�b�P���ȏ ����v���r����� :�(�^�����ğN��� ��ȯʯܯ� �6�x� ]���&���~�����Ŀ ƿؿ�P�5�t���h� Vό�zϰϞ����<� �L���@�.�d�R߈� v߬�����ߜ��� �<�*�`�N���߫� ��t���������8� &�\������L����� ��������4v�[ ��$�|���� �<!3��T �x����8 �,//</>/P/�/t/ �/��//�/?�/(? ?8?:?L?�?�/�?�/ r?�?�? O�?$OO4O �?�?�O�?ZO�O�O�O �O�O�O _bOG_�O_ z__�_�_�_�_�_�_ :_o^_�_Ro@ovodo �o�o�o�oo�o6o�o *N<r`�� �o����&�� J�8�n������^��� Z�ȏ���"��F��� m���6���������ğ ����`�E����x� f�������������8� �\��P�>�t�b��� ������$���4�ο(� �L�:�p�^ϔ�ֿ�� �����π���$��H� 6�l߮ϓ���\��ߴ� ������ ��D��k� ��4���������� ���^�C����v�d� ����������$�	 ������<r`�� ���� �$ &8n\���� ���/� /"/4/ j/��/�Z/�/�/�/ �/?�/?r/�/i?�/ B?�?�?�?�?�?�?O J?/On?�?bO�?rO�O �O�O�O�O"O_FO�O :_(_^_L_n_�_�_�_ �O�__�_o o6o$o ZoHojo�o�_�o�_�o �o�o�o2 V�o }�FhB��� 
��.�pU����� v��������Џ�H� -�l���`�N���r��� ����ޟ ��D�Ο8� &�\�J���n����� ݯ������4�"�X� F�|������l�ֿh� ����0��Tϖ�{� ��DϮϜ�������� ��,�n�Sߒ�߆�t� �ߘ��߼����F�+� j���^�L��p��� �����������$� Z�H�~�l�������� ������ VD z�����j��� �
R�y� B������/ Z�Q/�*/�/r/�/ �/�/�/�/2/?V/�/ J?�/Z?�?n?�?�?�? 
?�?.?�?"OOFO4O VO|OjO�O�?�OO�O �O�O__B_0_R_x_ �O�_�Oh_�_�_�_�_ oo>o�_eowo.oPo *o�o�o�o�o�oXo =|op^��� ���0�T�H� 6�l�Z�|�~���Ə� �,��� ��D�2�h� V�x�Ώ�ş����� ��
�@�.�d����� ʟT���P�ί���� �<�~�c���,����� ����ʿ�޿�V�;� z��n�\ϒπ϶Ϥ� ����.��R���F�4� j�Xߎ�|߲������� ���ߞ��B�0�f�T� ���߱���z������� ���>�,�b������ R������������� :|�a��*��� ����Bh9x lZ�~��� �>�2/�B/h/ V/�/z/�/��//�/ 
?�/.??>?d?R?�? �/�?�/x?�?�?O�? *OO:O`O�?�O�?PO �O�O�O�O_�O&_hO M____8__�_�_�_��_�_�_@_%od_nQ��$SERV_MA_IL  nUd`��JhOUTPUT�YhoP@�NdRV 2�V  g` (�Q4o�o�NdSAVEzlhiTOP10 2�i d j_ 2 DVhz���� ���
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�����U�eYP�oKcF�ZN_CFG �Ugc�d�a��eT�GRP 2�^��a ,B  � A��nQD;� �B���  B4~�cRB21�foHELLW��U��f�`�ou���%RSR��)�b� M���q�����ο��˿ ��(��L�7�pς�~���  �a�%�����Ϣ�����boP��������Ǌ��2oPd����ɦH�K 1׫  ߈߃ߕߧ������� ����%�7�`�[�m��������ìOM�M ׯ�ȢFTOV_ENBYd��a�iHOW_RE�G_UI7�LbIM�IOFWDL�x���l�WAIT4�A��v���t`X��d��TIMX������VAX`��l�_U�NIT3��iLC�Q�TRYX��e�N`MON_ALI_AS ?e��`heo�����
 t��#�GY k}�:���� ��/1/C/U/g// �/�/�/�/l/�/�/	? ?-?�/Q?c?u?�?�? D?�?�?�?�?O�?)O ;OMO_OqOO�O�O�O �OvO�O__%_7_�O [_m__�_�_N_�_�_ �_�_o�_3oEoWoio ozo�o�o�o�o�o�o /A�oew� ��X����� �=�O�a�s������ ��͏ߏ����'�9� K���o���������b� ۟������"�G�Y� k�}�(�����ůׯ� ����1�C�U� �y� ��������l����	� �ƿ?�Q�c�uχ�2� �Ͻ������Ϟ��)� ;�M�_�
߃ߕߧ߹� d�������%���I� [�m���<������ �����!�3�E�W�i� ���������n����� /��Sew�����$SMON�_DEFPROG &����� &*SYSTEM*��� 	�REC�ALL ?}�	� ( �}
xy�zrate 11� >192.16�8.1.15:16668 *=,�8 <Yk}�}!61A=O� �/� �./�g/ y/�/�0/�/T/�/�/ 	?/�/�/�/c?u?�? �/B?>?P?�?�?O�5�8copy fr�s:orderf�il.dat v�irt:\tmpback\�?�?hO�zO�O}/!Bmdb:*.*6OHOQO�O��O_�43x!D:\ �O+P�O�2�Oh_z_�_}4!Ua)_;_�?�_ �_o?(1�_�_�_ao so�o�?�?�?No�o�o o(?�o�o]o� �o�o8J��� $��Y�k�}��� 4�F�X������ ��� .�֏g�y�����0��� T����	��ğ��ҟ c�u�����B�>�P�� ���*���ί_�q� ������:�L�ݿ�� �&���ʿ[�m�ϒ� ��6�H��������"� ������i�{�ߠ�2� ��V������O0O�O �Oe�w��O7��OR� �����_-o?oP_a� s����_)�;������� �(��L�]o� ���A������ $���H�Yk}���� 3EX��� 2 ��g/y/�/�9/� T/�/�/	?��/R c?u?�?�+?=?��? �?O/*/�/N/_OqO �O�/�/CO�/�O�O_�X�$SNPX_�ASG 2����,Q�� P 0 '%R[1]@��,_WY?�C%W_�_ f_�_�_�_�_�_�_o �_7oo,omoPowo�o �o�o�o�o�o�o3 W:L�p�� ����� �'�S� 6�w�Z�l�������� Ə����=� �G�s� V���z���͟��ן� �'�
��]�@�g��� v��������Я��#� �G�*�<�}�`����� ��׿��̿���C� &�g�J�\ϝπϧ��� ��������-��7�c� F߇�j�|߽ߠ����� ������M�0�W�� f����������� ��7��,�m�P�w��� ������������3 W:L�p�� ���� 'S 6wZl���� �/��=/ /G/s/ V/�/z/�/�/�/�/? �/'?
??]?@?g?�? v?�?�?�?�?�?�?#O�DTPARAM �,U6Q W�	�'JP'D�@5'H~D�-PP�OFT_KB_CFG  fC2US�OPIN_SIM  ,[sF�O�O��Ov@=@RVNOR�DY_DO  �}E�ERQSTP/_DSB�NsBU_|aX=@SR �I� � &�@TY'LE1a_�\�T�C�TOP_ON_E�RR_;B�QPTN� �E�P��C�RRING_�PRM�_0RVCNT_GP 2�E:�A�@x 	Q_Po�h@>owobo�olWVD>%`RP 1LI�@�axI�g�o�o�o EBTfx�� �������,� >�P�b�t�������я Ώ�����(�:�L� ^�p���������ʟܟ � ��$�6�]�Z�l� ~�������Ưد��� #� �2�D�V�h�z��� ����¿����
�� .�@�R�d�vψϯϬ� ����������*�<� N�u�r߄ߖߨߺ��� ������;�8�J�\� n���������� ���"�4�F�X�j�|� �������������� 0BTf��� �����, SPbt����b�PRG_COUN�T�F��R�EN�Bo�M��D/_�UPD 1{[T  
�gBR/d/ v/�/�/�/�/�/�/�/ ?/?*?<?N?w?r?�? �?�?�?�?�?OOO &OOOJO\OnO�O�O�O �O�O�O�O�O'_"_4_ F_o_j_|_�_�_�_�_ �_�_�_ooGoBoTo fo�o�o�o�o�o�o�o �o,>gbt �������� �?�:�L�^������� ��Ϗʏ܏���$� 6�_�Z�l�~��������Ɵ�����_IN�FO 1@%s& H�	 ��c�N���r�?����@B�z=�����t���	�@���>�!�v�m�´�B������=�` @�� @���>��� >����� C�/�C�Q�Ch<C3����u��B������C�0B���Ã�G��Ҫ�9lw7��/��YSDEBU)G�A ��d))Q�SP_PASS��B?c�LOG �=�J!  r����  �%!��UD1:\x��#���_MPC���@%�#�@!̱A� �@!�SAV ����y���вC��׸SV�TEM_TIME 1���K  0  ¬�������ME?MBK  @%%!�����%�7�G�X;|& � @G���iߎߞ�b�����Y��^� y�@�� ��*�<�v�T�f�x�0������ ����� ��
��.�@�R�d�v��e������������ (:L^p� ������ ��SK�����@R�dX�� "�2(sߣ�p�� ��� ������%/7/I/[/O�u$� �u/��ߴ/`�/�/���/��?@'?9?K?]?o?�$s?�?���?�4^�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__�)�T1SVGUNwSPDy� 'c���4P2MODE_?LIM ��g�20T2=P]Q��/U�ASK_OPTI�ONX��g��Q_;DIr�ENB��5�c��QBC2_GRP 2#c����_̥"� C�c(\BC?CFG !�[~�� o"Ekem` eo���o�o�o�o�o�o �o?*cN` �������� �;�&�_�J���n�����ˏݏ�Ȍ��ɏ *�<����r�]����� ��H�ڟԯ����� ,��P�>�t�b����� ��ί������:� (�J�p�^��������� ܿʿ�� �6��� J�\�zόϞ���ϰ� �������.�@��d� R߈�v߬ߚ߼߾��� ���*��N�<�r�`� ������������ �$�&�8�n�\���H� ����������|�" 2XF|��n� ����0 fT�x���� �/�,//P/>/t/ b/�/�/�/�/�/�/�� 
??:?L?^?�/�?p? �?�?�?�?�? O�?$O OHO6OlOZO|O~O�O �O�O�O�O_�O2_ _ B_h_V_�_z_�_�_�_ �_�_�_�_.ooRo? jo|o�o�o�o<o�o�o �o<N`.� r������� &��J�8�n�\����� ��ȏ���ڏ���4� "�D�F�X���|���ho ʟܟ������B�0� R�x�f���������� ү���,��<�>�P� ��t�����ο���� �(��L�:�p�^ϔ� �ϤϦϸ������ȟ *�<�Z�l�~��Ϣߐ� ��������� ���D� 2�h�V��z���� ����
���.��R�@� b���v����������� ��N<r(� �����\��8&\Fz�$�TBCSG_GR�P 2"F��  �z 
 ?�  � �������5/�/Y/k+~�$�_d@ ��!?z	 HBLk(z�&~j$B$  C��0�/�(�/�/Cz�/(=�A�k(333?&�ff?��i%A���/m?80 k(�1͎6S5�0DHp?�=@�H0j%K1�5j$�1D"N!�?�?�?�?;O J�(I&�(nE�OLO^O �O�O�O�O�O_ [�H�:Q	V3.0�0�	lr2d S	*\PTTyk_f*_ �Q�I �Pt]�_  �_�_�[~J2�%�=Qo~�UCFG 'F�� �"j��Lb�R"owh�wo�o�jO�o�o�o �o�o=(aL ^������� ��9�$�]�H���l� ����ɏ��Ə���#� �G�Y��� d�v��� 2�����˟�ܟ� � 9�$�]�o�����N��� ��ۯƯ��zf6� BF�H�Z���~����� ؿƿ����2� �V� D�z�hϞόϮϰ��� �����
�@�.�d�R� tߚ߈߾߬����ߴ ����>�`�N��r� ����������&� ��6�8�J���n����� ����������"2 4F|j���� ���B0f T�x����� /�,//P/>/`/�/ 0�/�/�/l/�/�/? ??L?:?p?^?�?�? �?�?�?�?�?O O"O HOZOlO&O|O�O�O�O �O�O�O_�O_ _2_ h_V_�_z_�_�_�_�_ �_
o�_.ooRo@ovo do�o�o�o�o�o�o�o *�/BT� �������� 8�J�\��l������� ��ڏ����ʏ4�"� X�F�h���|�����֟ ğ���
���T�B� x�f���������Я�� ���>�,�b�P�r� t�����6Կ����� (��8�^�Lς�pϦ� �������� ߾�$�� H�6�X�~ߐߢ�\�n� �������� ��D�2� T�z�h�������� ������
�@�.�d�R� ��v����������� ��*N`
�x� �F���� $J8n��Pb ����/"/4/F/  /j/X/z/|/�/�/�/ �/�/?�/0??@?f? T?�?x?�?�?�?�?�? �?�?,OOPO>OtObO �O�O�O�O�O�Ol� _._�O_L_^_�_�_ �_�_�_�_ oo$o6o �_ZoHojolo~o�o�o �o�o�o�o2 V Dfhz���� ���
�,�R�@�v� d���������ΏЏ� ��<�*�`�N����� @_����ҟ|���&� �6�8�J���n����� ȯگ�����"��F��0�  l�p� �p���p��$TB�JOP_GRP �2(8���  ?�p�	�����*���@���@�� 0��  �� � � � ��p� @�l���	 �BL �  �Cр D�����<��E�A�S�<��B$�����@��?�33C�*���8œϞ�� �2�T�����;�2��t��@��?���zӌ�-�kA�>�Ⱥ�� �����l�>�~�a�s��;��pA�?��ff@&ff?�#ff�ϵ�8� ��L����}������:v,����?L~�}ѡ�D�H��5�;�M�@�33`�����>��|օ���8���`ự�	�D"��������`��r�|���"�9������g�v��x��� �������������� 0(V�b������p�C��p�	���	V3�.0�	lr2d��*b��k�p�{ E8� �EJ� E\� �En@ E��E��� E�� E��� E�� E��h E�H E��0 E� EϾ��� E���� E�x E��X F��D��  D�` E��P E�$��0�;�G�R��^p Ek�ui������(��� E�����?X 9�IR4! �H%�
z�`/r"�p�v#Ѭ߱/��E?STPARSI d�쵰��HR� ABL�E 1+��J p��(�' �k)�'��(�(o�w��'	��(
�(�(5p���(�(�(K!�#RDI�/��??(?:?L?^5�4O�?�;�? �?O O2N�"S�?�� �:�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo���@ �O��7�isO�O�O�O U?g?y?�?�?�8�"pb�NUM  8�U����x� J �K �"_CFG �,Y{s�@��IM?EBF_TT�!u8��� �vVERI#�az�v�sR 1-�+O 8mp�k�2� ;��o  �� �,�>�P�b�t����� ����Ώ�����(� :���^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�{�V�h� ��������¿Կ���H
��"�q_Sq�v@�u�� MI_CHA�N�w �u u�DB'GLV���u�u�!�x�ETHERADW ?�%���v ��������(x�R�OUT�p!WJ!�*�H��SNMA�SK���s��255.��N�ߖߨ�N�� OOLOFS_�DI� BŪ�OR�QCTRL .�{>Cw/&�T�J�\� n����������� ���"�4�F�X�j�z���������#PE_�DETAI����P�GL_CONFI�G 4Yyiq���/cell/$�CID$/grp1��;M_q�9C�߮���� �,>Pbt� �����/�� :/L/^/p/�/�/#/�/ �/�/�/ ??�/6?H? Z?l?~?�??1?�?�? �?�?O O�n}�?VO hOzO�O�O�Oq���O�M��?__1_C_U_ g_�?�_�_�_�_�_�_ t_	oo-o?oQocouo o�o�o�o�o�o�o�o );M_q � �������%� 7�I�[�m������� Ǐُ�����!�3�E� W�i�{������ß՟ ������/�A�S�e� w��������ѯ������ �Us�er View �)	}}1234567890J�\�n����������5�	̿��0�2=���� �2�@D�V�h�ǿٿ7�3� �����������o�1�߾4��j�|ߎߠ߲���#���߾5Y��0�B�T�f�x��ߙ�߾6 ���������,���M�߾7��������� ����?�߾8u�: L^p������� lCamera;�1� 0BT2BE�~ ��H�����//�  ���f/ x/�/�/�/�/g�/�/ ?S/,?>?P?b?t?�?�����?�?�?�? OO,O�/PObOtO�? �O�O�O�O�O�O�?�7 XىO>_P_b_t_�_�_ ?O�_�_�_+_oo(o :oLo^o_�72+�_�o �o�o�o�o�_*< N�or����� so���a�(�:�L� ^�p��������܏ � ��$�6���7t� ͏��������ʟܟ��  ��$�o�H�Z�l�~� ����I��7(	9�� � �$�6�H��l�~��� ۯ��ƿؿ���ϵ�ǧ9��O�a�sυϗ� ��P������Ϙ��'�@9�K�]�o߁�
	�0߼��������� ��:�L�^�߂��� ������ߕ�� ��� 5�G�Y�k�}���6�� ����"���1C U���I+����� �����1C� gy����h�� �;X//1/C/U/g/ �/�/�/��/�/�/ 	??-?��![�/y? �?�?�?�?�?z/�?	O Of??OQOcOuO�O�O @?��k0O�O�O	__ -_?_�?c_u_�_�O�_ �_�_�_�_o�O��{ �_Qocouo�o�o�oR_ �o�o�o>o);Mx_qm  i ���������0�B�T�f�    v~������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ�ؿj�  
`( � �p( 	 ���B�0�f�T� ��xϚϜϮ���������,���� � �oq߃ߕ������� ����c`�=�O�a� �߅��������&� ��'�n�K�]�o��� ������������4� #5GYk����� ����1 C�gy���� ���	/P-/?/Q/ �u/�/�/�/�/�// (/??)?p/M?_?q? �?�?�?�/�?�?�?6? O%O7OIO[OmO�?�O �O�O�?�O�O�O_!_ 3_zO�Oi_{_�_�O�_ �_�_�_�_oR_/oAo So�_wo�o�o�o�o�o o�o`o=Oa s���o�o��� 8�'�9�K�]�o�� �������ۏ���� #�5�|�Y�k�}�ď�����şן���B�"�@� �*�<�N���$����+frh�:\tpgl\r�obots\lr�m200id��_�mate_��.xml
���Ưد����� �2�D�V�F��� `���������Ϳ߿� ��'�9�K�b�\ρ� �ϥϷ���������� #�5�G�^�X�}ߏߡ� ������������1� C�Z�T�y������ ������	��-�?�V� P�u������������� ��);R�Lq ������� %7NHm� ������/!/�3/E.g��� |$�r�<< p� ?�E+�/E/�/�/ �/�/�/?�/?<?"? 4?V?�?j?�?�?�?�?��?�?�?
O8OF���$TPGL_OUTPUT 7P��P� h  tE�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo�'otEh �=@2345678901Lo ^opo�o�o�o�cF�Io �o�o�o/�o3@ew���Ez}� ����'���]� o���������O�ŏ� ���#�5�͏C�k�}� ������K�]����� �1�C�۟Q�y����� ����Y�ϯ��	��-� ?�ׯ�u��������� Ͽg�ݿ��)�;�M� �[σϕϧϹ���c� u���%�7�I�[��� iߑߣߵ�����q��߀�!�3�E�W���HA} c!�������������@j/�.�p* ( 	 1oc�Q��� u��������������� )M;q_�� �����7 %GI[��?f�f &��-�#/ 5//Y/k/9j��/�/ H/�/�/�/�/?,?�/ 0?b?�/N?�?�?�?�? �?>?�?O�?OLO^O 8O�O�O�?|O�O�OvO  __�O_H_�O�O~_ �_*_�_�_�_�_�_o l_2oDo�_0ozoTofo �o�o o�o�o�o�o. @dv�o^�� X����*��� `�r����������ޏ <�N��&���2�\�6� H��������ڟt�Ɵ �"���F�X���@��� (�z�į֯�����j� ��B�T��x���d��� ���0���Ϣ��>� �*�tφ�俪ϼ�Vπ��������(�:��)�WGL1.XM�L��o��$TPOFF_LIM �|���}��N_SV��  �����P_MON7 8������2y�STRT?CHK 9�������VTCOM�PAT��6��VW�VAR :��\Y�� � q�������_DE�FPROG %���%ZAD15 ADR*���z��_DISPLAY����ޡ�INST_�MSK  �� ���INUSER�,���LCK5���QUICKMENY����SCREx���7�tpsc@��5����ҩ�_���ST*��RACE_CFG ;���Y���	z�
?����HNL 2<��`� ��L^ p������
��ITEM 2=8� �%$12345678901  =<)Oai  !ow��3�z��A/ /w)/��v/��/ ��/�/M/=/O/a/{/ �/�/�/U?{?�?�/�? ?'?9?�?]?	O/OAO �?MO�?�?�?qO�O#O �O�OYO_}O�OX_�O s_�O�_�__�_1_�_ og_'o�_7o]ooo�_ {o�_	oo�o?o�o #�oG�o�o�oSk ��;�_q:� �U��y������� %��I�	�m��?�ŏ ��Ǐُ���w�!�͟ ��i�)�������+� ՟�������ůA�S� e��7���[�m�ѯy� ���п+��O��!� ��7ϩ�����߿��� ������K���oρϓ� ߷�c߉ߛ��Ͽ�#� 5�G�����}�=�O�� [����߲����1����g�����f���S���>k��  �k� ����
 ���������UD1:\&���}�R_GRP �1?� 	 @��q�m� ������� � �&J5nY?�  ����� ��/�//'/]/ K/�/o/�/�/�/�/�/��/	9�?%?{�S�CB 2@�� tq?�?�?�?�?�?��?�?Oq�UTOR?IAL A���LOv�V_CONFIG B�����	�O[MOUTPU�T C���@���O�O__1_C_ U_g_y_�_�_�_�_�_ �A�O�_oo1oCoUo goyo�o�o�o�o�o�_ �o	-?Qcu ������o�� �)�;�M�_�q����� ����ˏݏ���%� 7�I�[�m�������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ�������� '�9�K�]�o߁ߓߥ� �����������#�5� G�Y�k�}������ ����O�E�O'�9�K� ]�o������������� ������#5GYk }������� 1CUgy� ������	/ -/?/Q/c/u/�/�/�/ �/�/�/�/?/)?;? M?_?q?�?�?�?�?�? �?�?O?%O7OIO[O mOO�O�O�O�O�O�O �O_ O3_E_W_i_{_ �_�_�_�_�_�_�_o _/oAoSoeowo�o�o �o�o�o�o�oo+ =Oas���� �����&9�K� ]�o���������ɏۏ����������0�B�,��m���� ����ǟٟ����!� 3�E�W�i�������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sτ��ϩϻ������� ��'�9�K�]�o߀� �ߥ߷���������� #�5�G�Y�k�}�ߡ� ������������1� C�U�g�y�������� ������	-?Q cu������� �);M_q �������/ /%/7/I/[/m//� �/�/�/�/�/�/?!?�3?E?W?i?{?�;�$�TX_SCREE�N 1DD��,��}ip�nl/�0gen.htm�?�?�?OO�%O��Panel setup)L}�)OjO|O�O�O�O�OXONO�O__1_ C_U_�Oy_�O�_�_�_ �_�_�_n_�_-o?oQo couo�o�_,o"o�o�o �o)�oM�oq �����BT� �%�7�I�[�� �� ����Ǐُ���t�!� ��E�W�i�{��������>UALRM_M_SG ?�9��0 ���*��5�(� Y�L�}�p�������ׯ�ʯ����ӕSEV7  �Q�ђECFG F�5��1  �%@�  A��   ;Bȍ$
  ��# �5��ƿؿ���� ��2�D�V�h�v�]�GR�P 2Gg� 0��&	 ����ӐI�_BBL_NOT�E Hg�T��l�"�0�!�s���DEFPR�Oݐ%� (% �:ߖ (�a�L߅�p� �ߔ��߸������'���K���FKEYD?ATA 1I�9��Op v��&��������������,(��+��$(POINT  ]3�5����NCEL_����N?DIRECT����� EXT STE�P��6�TOUC�HU���ORE INFOO aH�l���� ��9 ]o� ��/fr�h/gui/wh�itehome.pngp��������point�*/</N/`/r/&�  FRH/FC�GTP/wzcancel/�/�/�/��/�/�#�indirec/4?F?X?j?8|?�/� nex#?�?��?�?�? O$�t?ouchup�?<O�NO`OrO�O$�arwrg�?�O�O�O �O_�8#_5_G_Y_k_ }_�__�_�_�_�_�_ o�_1oCoUogoyo�o o�o�o�o�o�o	 �o?Qcu��( �������;� M�_�q�������~�� ӏ���	��-�4�Q� c�u�������:�ϟ� ���)���;�_�q� ��������H�ݯ�� �%�7�Ư[�m���� ����D�ǿ����!� 3�E�Կi�{ύϟϱ� ��R�������/�A� ��S�w߉ߛ߭߿��� `�����+�=�O��� s�������\��� ��'�9�K�]����@����������v���������#5WiC, U�M����� �<N5rY� �����/�&/ /J/1/n/�/g/�/�/ �/�/���/?"?4?F? X?g�|?�?�?�?�?�? �?w?OO0OBOTOfO �?�O�O�O�O�O�OsO __,_>_P_b_t__ �_�_�_�_�_�_�_o (o:oLo^opo�_�o�o �o�o�o�o �o$6 HZl~��� ���� �2�D�V� h�z������ԏ� ��
���.�@�R�d�v� �������П���� ��/<�N�`�r����� ����̯ޯ���&� ��J�\�n�������3� ȿڿ����"ϱ�F� X�j�|ώϠϲ�A��� ������0߿�T�f� xߊߜ߮�=������� ��,�>���b�t�� ����K������� (�:���^�p������� ����Y��� $6 H��l~���� U�� 2DV�-�X�-�������}���,�/
/�/.// R/d/K/�/o/�/�/�/ �/�/??�/<?#?`? r?Y?�?}?�?�?�?�? �?O�?8OJO)�nO�O �O�O�O�O��O�O_ "_4_F_X_�O|_�_�_ �_�_�_e_�_oo0o BoTo�_xo�o�o�o�o �o�oso,>P b�o������ o��(�:�L�^�p� �������ʏ܏�}� �$�6�H�Z�l����� ����Ɵ؟����� � 2�D�V�h�z�	����� ¯ԯ������.�@� R�d�v���_O����п �����*�<�N�`� rτϖ�%Ϻ������� �ߣ�8�J�\�n߀� ��!߶���������� "��F�X�j�|��� /������������� B�T�f�x�������=� ������,��P bt���9�� �(:�^p ����G�� / /$/6/�Z/l/~/�/Т/�/�/���+�>������/? =�/7?I?#6,5Oz? -O�?�?�?�?�?�?�? O.OORO9OvO�OoO �O�O�O�O�O_�O*_ _N_`_G_�_k_�_�_ ���_�_oo&o8oG/ \ono�o�o�o�o�oWo �o�o"4F�oj |����S�� ��0�B�T��x��� ������ҏa����� ,�>�P�ߏt������� ��Ο��o���(�:� L�^�ퟂ�������ʯ ܯk� ��$�6�H�Z� l���������ƿؿ� y�� �2�D�V�h��� �Ϟϰ����������_ �.�@�R�d�v�}Ϛ� �߾���������*� <�N�`�r����� ���������&�8�J� \�n�����!������� ������4FXj |������ �BTfx� �+����// �>/P/b/t/�/�/�/ 9/�/�/�/??(?�/ L?^?p?�?�?�?5?�?��?�? OO$O6O��8K�����aOsO�M]O�O�O�F,�_�O�__�O2_D_ +_h_O_�_�_�_�_�_ �_�_�_oo@oRo9o vo]o�o�o�o�o�o�o �o*	�N`r� ���?����� &�8��\�n������� ��E�ڏ����"�4� ÏX�j�|�������ğ S������0�B�џ f�x���������O�� ����,�>�P�߯t� ��������ο]��� �(�:�L�ۿpςϔ� �ϸ�����k� ��$� 6�H�Z���~ߐߢߴ� ����g���� �2�D� V�h�?�������� ����
��.�@�R�d� v�������������� ��*<N`r ������� &8J\n�� ������"/4/ F/X/j/|/�//�/�/ �/�/�/?�/0?B?T? f?x?�??�?�?�?�? �?OO�?>OPObOtO �O�O'O�O�O�O�O_ _�O:_L_^_p_�_�_��_}��[�}�����_�_�]�_o)of,Zo~o eo�o�o�o�o�o�o �o2VhO�s �����
��.� @�'�d�K�����yﾏ Џ����'_<�N� `�r�������7�̟ޟ ���&���J�\�n� ������3�ȯگ��� �"�4�ïX�j�|��� ����A�ֿ����� 0Ͽ�T�f�xϊϜϮ� ��O�������,�>� ��b�t߆ߘߪ߼�K� ������(�:�L��� p�������Y���  ��$�6�H���l�~� ��������������  2DV]�z�� ����u
. @Rd����� ��q//*/</N/ `/r//�/�/�/�/�/ �//?&?8?J?\?n? �/�?�?�?�?�?�?�? �?"O4OFOXOjO|OO �O�O�O�O�O�O�O_ 0_B_T_f_x_�__�_ �_�_�_�_o�_,o>o Poboto�oo�o�o�o��o�o��{}������A@Se}=��sv,�� �}����$��H� /�l�~�e�����Ə؏ ����� �2��V�=� z�a�������ԟ���� 
���.�@�R�d�v��� �o����Я����� ��<�N�`�r�����%� ��̿޿��ϣ�8� J�\�nπϒϤ�3��� �������"߱�F�X� j�|ߎߠ�/������� ����0��T�f�x� ����=�������� �,���P�b�t����� ����K�����( :��^p���� G�� $6H �l~����� ��/ /2/D/V/� z/�/�/�/�/�/c/�/ 
??.?@?R?�/v?�? �?�?�?�?�?q?OO *O<ONO`O�?�O�O�O �O�O�OmO__&_8_ J_\_n_�O�_�_�_�_ �_�_{_o"o4oFoXo jo�_�o�o�o�o�o�o �o�o0BTfx ������� �,�>�P�b�t���]����]�����ÏՍ����	��,��:��^�E��� ��{�����ܟ�՟� ��6�H�/�l�S����� ��Ư���ѯ� �� D�+�h�z�Y����¿ Կ�����.�@�R� d�vψ�ϬϾ����� ��ߕ�*�<�N�`�r� ��ߨߺ�������� ��8�J�\�n��� !������������� 4�F�X�j�|�����/� ����������B Tfx��+�� ��,�Pb t���9��� //(/�L/^/p/�/ �/�/�/���/�/ ?? $?6?=/Z?l?~?�?�? �?�?U?�?�?O O2O DO�?hOzO�O�O�O�O QO�O�O
__._@_R_ �Ov_�_�_�_�_�___ �_oo*o<oNo�_ro �o�o�o�o�o�omo &8J\�o�� ����i��"� 4�F�X�j�������� ď֏�w���0�B� T�f�����������ҟh���� ���� ���!�3�E��g�y�S�,e���]� ί�����(��L� ^�E���i�������ܿ ÿ ����6��Z�A� ~ϐ�wϴϛ������/ � �2�D�V�h�w��� �߰��������߇�� .�@�R�d�v���� ����������*�<� N�`�r���������� ������&8J\ n������ ��4FXj| ������/ �0/B/T/f/x/�/�/ +/�/�/�/�/??�/ >?P?b?t?�?�?'?�? �?�?�?OO(O��LO ^OpO�O�O�O�?�O�O �O __$_6_�OZ_l_ ~_�_�_�_C_�_�_�_ o o2o�_Vohozo�o �o�o�oQo�o�o
 .@�odv��� �M����*�<� N��r���������̏ [�����&�8�J�ُ n���������ȟڟi� ���"�4�F�X��|� ������į֯e������0�B�T�f��$U�I_INUSER  �������  �g�k�_MENH�IST 1J���  (� ����*/S�OFTPART/�GENLINK?�current=�editpage�,ZAD15,1 ���-�?��(���menu��153 ϛϭϿ����߿��1��!�3�E�W������2ߥ߷����� j�|��(�:�L�^������4�����&��'t�v�2�-��?�Q�c�^����48�,2h������������۱��
.@Rdv ��� ����+=O as����� �/�'/9/K/]/o/ �//�/�/�/�/�/�/ �/#?5?G?Y?k?}?�? ?�?�?�?�?�?O�� 1OCOUOgOyO�O�O�? �O�O�O�O	__�O?_ Q_c_u_�_�_(_�_�_ �_�_oo)o�_Mo_o qo�o�o�o6o�o�o�o %�oI[m ���D���� !�3�O<�i�{����� ��Ï������/� A�Џe�w��������� N�П����+�=�O� ޟs���������ͯ\� ���'�9�K�گ\� ��������ɿۿj��� �#�5�G�Y�D��� �ϳ���������� 1�C�U�g��ϋߝ߯� �������߆��-�?� Q�c�u������� ������)�;�M�_� q�������������� ��%7I[m�j��$UI_PA�NEDATA 1�L�����  	�}�/frh/gu�i�dev0.s�tm ?_wid�th=0&_height=10� �� ice=TP&�_lines=1�5&_colum�ns=4� fon�t=24&_pa�ge=whole�� �h�)pri9m/X  }[`����� )� ��#/
/G/Y/@/}/ d/�/�/�/�/�/�/?��/1?h��� �    ][�in?�?�?�? �?�??�?_O"O4O FOXOjO�?�O�O�O�O �O�O�O�O__B_T_ ;_x___�_�_�_�_E7 � �U�Oo$o6o HoZolo�_�oO�o�o �o�o�ouo2D+ hO������ �
���@�'�d�v� �_�_����Џ��� Y�*��oN�`�r����� ����!�ޟş��&� 8��\�C�����y��� ��گ�ӯ�����F� X�j�|������Ŀֿ I�����0�B�Tϻ� x�_ϜϮϕ��Ϲ��� ���,��P�b�I߆� mߪ��/������ (�:�L��p�㿔�� ��������U��$�� H�/�l�~�e������� �������� DV ���ߌ����� 9
}�.@Rdv ������/ /�</#/`/r/Y/�/ }/�/�/�/�/cu&? 8?J?\?n?�?�/�?�? )�?�?�?O"O4O�? XO?O|O�OuO�O�O�O �O�O_�O0_B_)_f_0M_�_�/?}��_�_ �_�_
oo.o)�_So �5Boo�o�o�o�o�o @o�o�o!W> {b���������/��83;�$�UI_POSTY�PE  5� 	 ;����a�QUICKM_EN  p�����c�RESTOR�E 1M5�  ��*default��;SINGL�EԍPRIM�ԏmmenup�age,148,2 1<�q������� J���П������� <�N�`�r����"��� ���ϯ��
��.�@� �d�v�������O�п �����ï%�7�I� ���ϖϨϺ���o��� ��&�8�J���n߀� �ߤ߶�a�������Y� "�4�F�X�j���� ������y�����0� B�����a�s������ ��������,>P bt�����ޚ�SCRE��?���u1sc��u2!3!4�!5!6!7!8�!�TATl�� �ă5Y�USER�ks#�3��4�5�6�7�8�a�NDO_?CFG Np��P��Qa�OP_CRM�5  �U&a�P�Dd���None���_I�NFO 1O5f 0%��/�8 o/�/�/�/�/�/
?? �/@?#?d?v?Y?�?�?��?�?��S!OFFS�ET Rp�j! �?����!O3OEOWO �O{O�O�O�O�OO�O ___J_A_S_�_w_��_�_�Kŏ�]�_
o
��_/o�8UFRAM�%�/P!RTOL_�ABRTSoN#kbE�NBtoehGRP �1S����Cz  A��c�a��o�o�o�o"v,>cj⯀U�h#!�kMSKG  �ef!�kNPa%^)�%�_��eO_EVNs`�t&��v�2T�;
 h�#!UEVs`!�td:\eve�nt_user\��7�C7<�o� F�q�/�SP5�:�spotweldl�!C6��r���#�t!�K�	�>��q ��-��q���Q�c�ܟ �� �����ϟH��l� �)�_�����د���� ˯ ��D���z�%� ����[�m�濑�
ϵ��Ǻ�WRK 2U��a8�nπ�  \ϥϷϒ�������� #���G�Y�4�}ߏ�j� ���ߠ��������1���B�g�y��$VA�RS_CONFI��V�; FP�݈��CMR�b2\N�;xy� 	$ ���01: SC�130EF2 *(�	����X�ȸpm�  #!?�p�@pp"p�z� 	o]�g���������������`�uA�����,� B���G�K ��l���_��� ����2�h�Se�Q����IoA_WOF�]^-˶,		�Q;%/>+'G�P �> ����RTWINUR�L ?�������/�/�/�/�/�/��SIONTMO�U� ��%��^S۳�S۵�@�a FR:}\�#\DATA؏�  �� U�D166LOGC? � \9EXh?'q'� B@ ���2{1U��?{1�?�?�θ � n6  ������2zt��`F��  =���BA��?@|=TRAIN�?AQB�d�CpBEFF/B�0�(��_� ( ��I�M��O�O�O_ _P_>_t_b_|_�_�_p�_�_�_�(_GE3`�/C�
�`'p4b,
g�0RE!0a�i��.��LEXdb�����1-e�/VMPH?ASE  ����C ��RTD_F�ILTER 2c.� �&��T��o +=Oas� ����o�������1�C�U�g��)SH�IFTMENU {1d�K
 <�<1%�?ŏ2����ɏ �ُ�8��!�n�E� W�}��������ß՟�"���	LIVE�/SNA��%v�sfliv�n4����# SETU<��W�menum�r�@�ѯ�"��3e`+�|�MO3ftn�z���ZD�gQm˳<��A�P�$WAITDINEND8�L!�k�OK  ��醼 :��S����T�IM5���G r�͔�%˴��ӿ�<򿆸RELE�a5���k��/6m�_AC�TJ�4� !��_?1 h��%�5߅���RDIS�����$XVRnai~tn�$ZABC��;1jQk ,�@��2=��-ZIP2kQo���)����MPCF_G 1	l��l!0L"��q�7�MP��m����P���c���`�*�  6n�G�6��"IG�o�5�j�5�i���A�H�C�/��CQ�Ch<��0�Q���;=��/";��P������ɿN?���������������6�?6��lT����@�?���,������p9�������C�C��0B��Ã��G�Ҫ�9l�w7³��,�I�䮵9lfw$@�PJ\�r��������6 �����J�p`n��_CYLIND�a�oR� �p6 ,(  *o�w3`l���� �� //'.iJ/�n/U/ g/�/��/�/�///? �/�/F?-?j?Q?�/�?Ȳ?�Cp*� �g��?L^���6O!O�ZO?I�?�O?G��AA��=SPHERE 2qO�?�OT? �O_�O:_�?�Op_�_ �/�_E_+_�_�_ o�_ Y_6oHo�_�_~o�_�o �o�o�oo�o ��ZZ�� ��