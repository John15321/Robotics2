��   ��A��*SYST�EM*��V9.1�0185 12�/11/2019� A 
  ����DRYRU�N_T  4� $'ENB � $NUM_�PORTA ES�U@$STAT�E P TCOLu_��PMPMCm�GRP_MASK�ZE� OTION�NLOG_INF�ONiAVcFL�TR_EMPTY�d $PROD_�_ L �ESTOP�_DSBLAPOW_RECOVA�OPR�SAW_�� G %$I�NIT	RESUME_TYPEN�DIST_DIF}FA $ORN4�1� d =R���&J_  4� $(F3ID1X��_ICIf�MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�� �MKR-�  $LIN�c   "_S�IZc�� �. �X $USE_FLC 3!�:&iF*SIMA7#Q�C#QBn'SCAN��AX�+IN�*I���_COUNrR�O( ��!_TMR�_VA�g# h>�ia �'` ����1�+WAR��$�H�!�#Nf3CH�PE�$,O�!PR�'Ioq6��OoATH-� P $ENA#BL+�0B�T���$$CLA�SS  �����1��5��5�0V�ERS��7�  �iAIRTU� �?@'/ �0E5���"����@kF1@�1pE��%�1�O���O�Ob����AEI2LK �O+_=_O_a_ s_�_�_�_�_�_�_�_�oo'o9o�O)W?yHW@ �� zj�0�o�o�i�� �� 2LI  #4%Ho�o��mA}A �o+
Oa@�� v������'� ��]�<�}A�c$"+ (�k�K@����pA��X��0A@�N� ����0�B�T�f�x� ����������pF}AՁ }A����*�<�N�`� r���������̯ޯ�4rhM��C� 2�lՏ;�M�_�q��� ������˿ݿ��� Ԝ-�F�X�j�|ώϠ� ������������)� B�T�f�xߊߜ߮��� ��������,�7�P� b�t��������� ����(�3�E�^�p� ��������������  $6A�Zl~� ������  2DOhz��� ����
//./@/ K]v/�/�/�/�/�/ �/�/??*?<?N?Qh �4�0���?=@