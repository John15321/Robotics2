��   ��A��*SYST�EM*��V9.1�035 7/1�9/2017 �A   ����BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG����DHCP_CTR�L.  0 �7 ABLE? $�IPUS�RET�RAT�$SE�THOST��N�SS* 8�D��FACE_NU�M? $DBG_�LEVEL�OMo_NAM� !� {FT� @� �LOG_8	,CM�O>$DNLD_FILTER��SUBDIRCA�PC��8 . �4� H{ADD�RTYP�H N�GTH�����z +LSq D� $ROBOTyIG �PEER�ބ MASK�MR�U~OMGDEV�����PINFO~�  $�$$TI ���RCM+�8 ?$( /�Q�SIZ�!S� T�ATUS_%$MAILSERV� $PLAN� �<$LIN<$�CLU��<$T�O�P$CC�&F�R�&YJEC|!�Z%ENB � A�LAR:!B�TP�,�#,V8 S���$VAR�)M�O�N�&���&APPL��&PA� �%��'P�OR�Y#_�!�"A�LERT�&i2UR�L }Z3AT�TAC��0ERR�_THROU3US0�9H!�8� CH- c%�4MAX?WS_�|1��1MOD��1I�  �1o }(�1PWD  � cLA��0�ND�1�TRYFDELA�-C�0G'AERSI���1Q'ROBICL�K_HM 0Q'� XM�L+ 3SGFRM2U3T� !OUU3 3G_�-COP1�F�33�AQ'C[2�%�B_AU�� 9 R�!�UPDb&PCOU�{!�CFO 2 
$V*W�@c%�DUMMY1TW2^?�RDM* �$DIS��S)N,#	3 �	o!��"%"_WI�CT?Z_INDE�3�PgOFF� ~UR�Y�D��S�  
o t Z!RT�0�N�cD�bHOUU#E%Af:a"f:a�1fLOCA� #{$NS0H_HE�K��@I�/ 3 �$ARPH&�_7IPF�W_* O2�F�PQFAsD90�VHO_� 5R{b;EL� P��r�90WORA�$ACCE� L�VO#�FS1�IcCE�3p� �$�c  ���RqJ��
��
Gp�PS�A�Pw# ��cqIz0ALOaq'�0 px
���F��p��{p�r�u�$� 2�{ "��]r@�}�p�� �}��!Yq�A����$� _FL�TR  oy�p U��������U��$�}2U��bSH[AR� 1�y P=���t��� C��g�*���N���r� ��埨�	�̟-��Q� �u�8�J���n�ϯ�� 󯶯�گ�M��q� 4���X���|����޿ �ֿ7���[��g�B� �ϵ�x��Ϝ�����!� ��E���{�>ߟ�b� �߆��ߪ߼����A� �e�(��L����`����Y�z _LUA�1n�x!1."B�0���A�1R���255.��I�����u@�2G�Y��� m��������3��Y�@6 ����	��47�Y�� ]o����5 �Y�&�����6'Y��M_q����7!"�S���S��܀ �� Q� ���<9/n/�/ S/�/�/�/�/�/�/��P�/.?@?R??v?�?��?�?k?�?�?�?���?���u>O)L
Z�DT Statu�s�?MO�O�O�O��}�iRConnect: irc�D//alertkN �O_"_4_�G}Ob_t_��_�_�_�_���sP�"��d���_�_	o o-o?oQocouo�o�o�o�o�o�s$$c9�62b37a-1�ac0-eb2a�-f1c7-8c�6eb56b02a8  (Q_"uO FXj|�����((�0"�r2J�u 0�v3C5 �,$=� ��3��%��I�0�V� �f�����Ǐُ���� �!���W�>�{�b����0!/� DM_�!/��SNT-P��	��%u��������������#ϓUSTOM' 
�����/ � ��$TCPIP����0H'%!�TEL'�/�,!��H!T�R�����rj3_tp�d)O 4��!KCLƯ˫���v!CRT%��l��'"��!CON�Sm�̪ڡib_Osmonu�i�