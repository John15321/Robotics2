��   K�A��*SYST�EM*��V9.1�035 7/1�9/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_���$$C�LASS  ������D��D�VERSION�  ���/IRTUA�L-9LOOR� G��DD<x$?������kn,  1 <DwX< y�����C�����	/��Z�Zm//�/_/p�/�/�/$ �/��/	?';�$MNU�>A\"�  <������3��g0��6 �"!�ik0�4x0s1D��B� �zP%��?��?�? �?�?�?OOOQO7O IOkO�OO�O�O�O�O�_�O�O_M_�;5N_UM  �����w92TOOLC?�\ 
Y;)-4���5���PSQ,�V�a�kBCv�7_Y_	o1_o?o%o 7oYo�omo�o�o�o�o �o�o�o;!Cq Wy�����sV �Q�Vy�[