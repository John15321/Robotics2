��   ?Q�A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����MN_MC�R_TABLE �  � $M�ACRO_NAM�E %$PR�OG@EPT_I�NDEX  �$OPEN_ID�aASSIGN_7TYPD  qk�$MON_NO�}PREV_SU�By a $USE?R_WORK���_L� MS�*RTN  �&�SOP_T � � $�EM�GO��RES;ET�MOT|�GHOLl��1�2�STAR PGDI8G IAG�BGC�TPDSN�REL�&U�� �� �EST����SFSP�C���C�C&�NB��S)*$T8*$3%)4%)5%)�6%)7%)S�PN'STRz�"D�  ��$$CLr   �����!������ VERSI�ON�( � �i�!IRT�UAL�/�!;LDUIMT  ���� ���4MAOXDRI� ��5�
4.1 �%� � d%�Open ha�nd 1����%� ?�? �"  �13�0ClosAeo?�?�?	O�9�7Relax�?�?GO$mO�9�6j82oOPO�OtO�3�?�O�O&_ �O�6 +O__�_;_�4�F�_�_�_�_�[ �3��(@�_6o�_Zo	o o�o?o�o�ouo�o�o �o �o�oVS� ;M�q���� .��R�����7��� [�m����ߏ�Ǐُ N���r�!�3�m���i� ޟ�����ß8�J��� 3���/���S�e�گ�� ׯ���ѯF���j�� +�������ֿ����� ��0�߿�+�x�cϜ� K�]��ρ��ϥϷ��� >���b��#ߘ�G߼� ��}߷���(����� ^��[��C�U���y� ����$�6�!�Z�	� ���?���c�u����� �� ����Vz) ;u�q��� �@R;�7� [m���/�� N/�r/!/3/�/�/�/ �/�/�/?�/8?�/�/ 3?�?k?�?S?e?�?�? �?�?�?�?FO�?jOO +O�OOO�O�O�O�O_ �O0_�O�Of__c_�_ K_]_�_�_�_�_�_,o >o)oboo#o�oGo�o ko}o�o�o(�o�o ^�1C}�y ���$��H�Z�	� C���?���c�u�ꏙ� � �Ϗ�V��z�)� ;�����柕���� ˟@���;���s��� [�m�⯑����ǯ� N���r�!�3���W�̿ ޿��ǿ�ÿ8���� n��kϤ�S�e��ω� �ϭϿ�4�F�1�j�� +ߠ�O���s߅߿�� ��0�����f���9� K���������,� ��P�b��K���G��� k�}�������(���� ^�1C��� ���$�H�	 C�{�cu�� /��	/V//z/)/ ;/�/_/�/�/�/�/? �/@?�/?v?%?s?�? [?m?�?�?O�?�?<O NO9OrO!O3O�OWO�O {O�O�O_�O8_�O�O n__�_A_S_�_�_�_ �_�_�_4o�_Xojoo So�oOo�oso�o�o�o �o0�o�of�9 K������,� �P���K������� k�}�򏡏�ŏ׏� ^����1�C���g�ܟ �ן$�ӟH���	� ~�-�{���c�u�ꯙ� ���ϯD�V�A�z�)� ;���_�Կ����Ͽ� �@���v�%Ϛ�I� [ϕ��ϑ�ߵ���<����`�r�!�[�
Se�nd Event�s�S�SENDEgVNT��Q�և�� %	��Datya�߶�DATA�������%��Sy�sVar;��SY�SVw����O�%�Get�x�GE�T+��޳�%R�equest M�enu���REQOMENU?����� ]ߞ�Y���}�+����� .��d�7 I�m����* �N����� i{��/��/ \/G/�///A/�/e/�/ �/�/�/"?�/F?�/? |?+?�?�?a?�?�?�? O�?�?BO�??OxO'O 9O�O]O�O�O�O__ _>_�O�Ot_#_�_G_ Y_�_�_�_o�_�_:o �_^oooYo�oUo�o yo�o �o$6�o l�?Q�u� ���2��V��� ������q������� �ˏݏ�d�O���7� I���m�⟑���ݟ*� ٟN������3����� i���𯟯�ïկJ� ��G���/�A���e�ڿ �����"��F���� |�+Ϡ�O�aϛ����� ߻���B���f��'��a߮�]��߁ߓ��$�MACRO_MA�XX�������Ж�SOP�ENBL ���2��ݐѐ��_���"�PDIMS�K�2�<�w�S�U���TPDSB�EX  K��U)�2�����-�