��   v��A��*SYST�EM*��V9.1�035 7/1�9/2017 �A   ����UI_CONF�IG_T  �X J$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY7]0�ODE�
1CWFOCA �2C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_Gv!k FKE�E ��3;CSP_NAM��#DIMC4:1YABRIGH83s kDJ7�CH91&USTO�[@  t v@AR$@PIDDr�BC�D*PAG� �?dAEVICE��ISCREuEF����GN�@$FwLAG�@��&��1  h 	$�PWD_ACCE	S� =E8�HS�:1�%)$LABE�� $Tz j�(P�3vR�	SUS�RVI 1  < `kR*kR�lQ7PRI�m� t1��PTRIP�"m��$$CLA3P O����Q��R��R�P\ SI��W�  ���QIRTs1�_�P'�2 L1W�L1a��R	� ,��$?���_b`hcdc�^a�� , ��  �o��
 ���Q�o�o�o�o#5 �oZl~ ���C����  �2��V�h�z����� ��Q����
��.� @�Ϗd�v��������� M������*�<�N� ݟr���������̯[� ���&�8�J�ٯn����������ȿڿ_`?TPTX����j�	�� s ��綄�$/sof�tpart/ge�nlink?he�lp=/md/t�pmenu.dg@ܿvψϚϬ�e�&A�S�pwdb����� /�d�S�e�w߉ߛ߭� <���������+�� ��a�s�������+��Q�f�fbc��($P������4��X����Qba~�o赊�~�|�L���c���aH���H��H�  H�	F��K����淤��`���`  ���F QO���I#H�qFG�8c�B 1	h�R \��_��� RE�G VED=����wholemod�.htm�	sin�gl�doub~�tripbrows) `�_q�M�� ���/����_dev.s�le/4} 1h,	t�/7 }//A/�/�/?�/+?�=?O?a?s?�?�  (`�?�?�?�?�?O O02ODOVO`F @�?�O �OfO�O�O�O�F�	�? �?_%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWo%'ooio�o �o�o�o�o�o' 9K]o���� ���?�(�:�L�^� p����������O܏� ��Ϗ$�6��O�O�~� y�����Ɵ��ӟ�� 	��-�V�Q�c�u��� ����yo˯ů��� )�;�M�_�q������� ��˿ݿ���%�7� �rτϖϨϺ����� �����8�J��+� �ߒ�I�[�A������� ��"��/�A�j�e�w� ������������ կ'�!�O�a�s����� ����������' 9K]o��a�� ��(:L^ pkߔ�u��� �߷ߝ6/1/C/U/~/ y/�/�/�/�/�/�/? 	??-?V?Q?c?1��? }?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O�*_<_N_ `_r_�_�_�_�_�_���_o�_�_8oJoXj��$UI_TOPMENU 1#`�yaR 
�d{aQ)*d?efault_�M�*level�0 *�K	 ��o�0�o�o�o�btpio[23]�8tpst[13x�O�o�o�=h�58E01_l.�png��6me�nu5�y�p�q13�z�r�z�t4�{��q��5�\�n������� ��RJ�ߏ���'��9�Ȅprim=��qpage,1422,1@�y����� ����̏���	��-��?�ΖT�class,5H�}�������4ůД\�13̯���&�8�J�ѓT�53f���������οѓT�8u�	��-�?� Q�ПuχϙϫϽ����I|`ya�o߶m��`�q��1�O�9vtyD}<,>qmf[0FD�}	|�c[1643w��593x�q�e���x2��}G��z	��w �{��E���������� ��e�>�P�b�t��� ��'�����������[�2(]o�� �4f����# ���dv���[�m�1����/ /�2/��T�ainedi��i/{/�/�/�/���config�=single&>T�wintp`��/ �/? ?2?�J{a��@? l?�et?��?�?�? �?�?OO'O�?3O]O pO�O�O�O�O�O�O9� �O$_6_H_Z_l_~_�� �_�_�_�_�_�_�_ o 2oDoVohozo	o�o�o �o�o�o�o
�o.@ Rdv���� �����<�N�`� r�����%���̏ޏ�� ����8�J�\�n������N��ȟ�%�K;��O���s�0�U���=�u�����d�b��(��L���B�0�6=�u7u���� ��˿ݿ(���%�7� I�[��ϑϣϵ���(�����"�1�%� 7�I�[�m�xϑߣߵ� ������z��!�3�E� W�i�{�|������������6 �5�G�`Y�k�}��$w�74�� ��������L<��4�5	TPTX[2c09��TDO24��0"�|Z�O18t�P��Wj0�2��`WA���3��tv8��*<N$0f#1�f_�S:�$tre�eview�#}�3���&dual=o��81,26,4 �'/9/K/
�o/�/�/ �/�/�/X/�/�/?#?�5?G?��;�z�53 �$���?�?�?�/�? OO1OCOUO�?yO�O��O�O�O�OZ?l?��1��?$2�>_P_b_ �6�O��edit ��_(_�_�_�_��� ���_�S�_GoYoko lo�o㕠o�o��o �o'9Kp�o i������ � �o�)�P�b�t����� ��iOΏ�����(� ��L�^�p�������5� ��ܟ� ��$�6�ş Z�l�~�������C�د ���� �2���D�h� z�������¿Q���� 
��.�@�Ͽd�vψ� �ϬϾ�moo�ϣo� �;�M�_�q߄ߕ� �߹�'�������%� 7�I�[�m�/������ �������[�4�F�X� j�|������������ ����0BTfx ��+���� �>Pbt�� '����//(/ �L/^/p/�/�/�/5/ �/�/�/ ??$?���� Z?	�~?�߃�?�?�? �?�?�?OO�?+OUO gOyO�O�O�O�O�O�� 
__._@_R_d_v_�/ �_�_�_�_�_�_�_o *o<oNo`oroo�o�o �o�o�o�o�o&8 J\n���� ����"�4�F�X� j�|������ď֏� �����0�B�T�f�x� ��9?K?��o?�KO�O ��+�=�O�a�t��� 󟑯��ͯ߯��� '�9��Op��������� ʿ�ܿ ��$�6�H� Z��~ϐϢϴ����� g���� �2�D�V��� hߌߞ߰�������u� 
��.�@�R�d��߈� ��������q���� *�<�N�`�r�������������������*default���Ξ*level�8W���O�m �tpst[1�]{	�y�tpio[23����u�Z�"4m�enu7_l.pkng7T13YBf5nS�Q4�u6Yf����/ #/5/��Y/k/}/�/�/ �/B/�/�/�/??1?�C?�"prim=�Tpage,74,1H??�?�?�?�?��"\6class,13�?OO&O8OJO�?�25PO�O�O�O�O�O�#�<tO__`,_>_P_S?e218l?��_�_�_�_�_�O�26��_o#o5oGoYo8��$UI_USERVIEW 1�����R 
��`oڒ�o�o3m�o�o�o#5 �oYk}��D� �����o�,�>� �y���������d�� ��	��-�?��c�u� ������V���ʟܟN� �)�;�M�_������ ����˯n����%� 7���V�h�گ���� ǿٿ�����!�3�E� W�i�ύϟϱ����� �������x�A�S�e� w߉�,߭߿������� ��+�=�O�a�s�� ����������� '���K�]�o�����6� ������������� 0��T}���� h��1�U gy��H��� @	//-/?/Q/�u/ �/�/�/�/�/r/�/? ?)?;?�H?Z?l?�/ �?�?�?�?�?�?O%O 7OIO[O�?O�O�O�O �Or?|O�O�OjO_E_ W_i_{_�_0_�_�_�_ �_�_�_o/oAoSoeo h