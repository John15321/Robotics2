��  	w^�A��*SYST�EM*��V9.1�0185 12�/11/2019� A  �����AAVM_�WRK_T  �� $EXP�OSURE  �$CAMCLB�DAT@ $PS_TRGVT��$X aH]ZgDISfWg�PgRgLENS_CENT_X��YgyORf  � $CMP_G�C_�UTNUM�APRE_MASwT_C� 	��GRV_M{$�NEW��	ST�AT_RUNAR�ES_ER�VTSCP6� aTCb32:dXSM�p&&�#END!�ORGBK!SMp��3!UPD�O�ABS; � P/ �  $P�ARA�  ����AIO_wCNV� l� �RAC�LO�M�OD_TYP@F+IR�HAL�>#�IN_OU�FA�C� gINTER�CEPfBI�I�Z@!LRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CESI0�!H1�!"PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W� @V�R!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2 � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1 UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t�cbMO� �sE 	� [M�s��2�wREV�BILF��!XI� %�R 7 � OD}`j��$NO`MD�+� `�x�/�"�u�� ����^��@D�d p E R�D_Eb��$F�SSB�&W`KBD�_SE2uAG� G
�2 "_��B�� V�t:5`ׁQC���a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR��BIGALLOW� (KD2�2�@VAR5�d!�A>B ��BL[@S � ,KJqM�H`9S�pZ@M_O]z�ޗ�CFd �X�0GR@��M�NFLI���;@UIRE�84�"� �SWIT=$/0_N�o`S�"CF_�G�� �0WAR�NMxp�d�%`LI��V`NST� CO�R-rFLTR^�TRAT T�`>� $ACCqS��� X�r$ORIأ.&ӧRT�`_SYFg��HGV0I�Ep�T��PA�I��5T���HK�� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8�  �0��x@�2� @� TRQB��$%f��ր����c_U���� COc <� ����Ȩx3�2��LLECM�}-�MULTIV4��"$��A
2FS�I�LDD��c� DET}_1b  4� STY2�b4�=@��)24��e`DԼ� |9$��.p��6�aI`�* \�TO�:�E��EXT����p���B�ў22�0,D��@��1b�.'�B ��G�Q� �"Q�/%�a��X� %�?sdaD�U� Sҟ؈;A�Ɨ�M�� �� CՋO�! L@�0a�� X׻pAβ$JOBB���֍�v��IGO�" dӀ �����X�-'x���G��ҧ]�C�`��b# etӀF� �CNG�AiBA� ϑ��!��� /1��À�0����R0aP/p3���$
��|��BqF]�
2J�]�_RN��C`J�`�e�J?�D/5C��	�ӧ��@����Pr�O3л!% \�0�RO�6� �IT<�s� NOM_8pn#��c ���TU��@P� � ��&"+P��� ӨP�	ݭ��RAx@n �3�A����
$TF3%#D%3
T��wpU�13��}�%mHrzT1�E���ޣ�#ݤp�%ߢQlYNT�"�� DBGDE�!'D�]�PU���@t����"��AX��"�uwTAI2sBUFۆ;%�1( ��P&V`[PI84'mP�'EM�(M�)B �&F�'�SIMQS�@ZK;EE3PAT�z�`�8"�"�MC��1)S�0��`JB�����aDECg:� g5e������* �U�CH�NS_EMPͲ#$G��7�_��c�;�1_FP)�TC�6S���5�`%��4�} ��V����W���JR����SEGF�RAq�O�� #PT�_LIN�KCPVAF���`  C$+�� �ckBZ��PBzr���@>6,` +�Ԧ ��A�0��Ad0o`Arp�D���Id1SIZh���	T�FT�C�Z1Y�ARSm��CP@'�@Ic\1@cX�0<@L��8��0�VCRCߥ�sCC���U1@�X�1��2�Mpq�U�1`�XD�Q�UDݤأiCk �p��
DK`݀f��RhSEVRf �Fha_	EF�0N�f�Pd1�&hB��5�jC}�+�OVSCA[��A�f����13��-�	<�ׇMARG���"a�F@@���1DcQ�rN�0LEW�-��R��P<��o�l��RɄ.� ����ǯ��� 5ڡR�`HANC��$LG5��a��Ӑ��ـF��Ae����0RYr�3
����
��@ �RA��
�AZ��0Q�N`�O��FCT��sp�F��R�0\P0b ADI��O�� +���+���&���5�5Є���S[�g���BMPUD(PY�1��GAESCPjc��W��%N  S-��U0ۑuU�/)�TIT'q�<�b�%ECA:!�!E'RRLd��0�&Q��OR�B$������~Ұ$RUN_O��SYS��4������u�REV�V@��?DBPXWO�P�=10�$SKo�"�1�DBT�pTRLn�2 �C AC��0��%�m�U DJ�p��_�`�!A�ǀM�P5L�A_2WA��j�EE��D!w�!%R|hO�UMMY9��ڠ�1� ��DBd[��3���!PR�Q� 
��ٱ9��4� г$r��$ Q��Lة5L�z����6�^z�PC�7*��<�ENEC0Tq�8I�����RECO}R$�9H mގ�4$L��5$ أ�"E���R@��VA��s_Dց� ROS �"SK�����I�=�א��PA��JVB�ETURN���SMeR(�U #�CRʰ�EWMDB0GNsALV �"$LA� �[�*6$P-�g7$Pv�s�8o��!�PC��#�DO�^@-�Ŵ���R˶GOg_AW�ܱMOz���p���CSS_+CN4�YO�:��T���0���ID�T�2*��2�N��O@�J���v`Iְ ; oP $>�RB�B���PI�POl�IG_BY��vЅ�TVR���HNDG$�< H�`�1a�@cS��DSBLI��s��ְ0}����LS$�=0��0� ��FB�FEձL�9����5z��>D�$DO�1�C�pMC�0q��4(��9�RH��W��K�4ELE�ur�
^��SLAVr?xB�INS ���#����_R@P�@\`�pS� }�l�}�l�{u��[!e��ے�I���B�r�W��D�NTV�#��VE�$��SKI lA4;3��2UB�1�J�f�1C�
DSAF�7�5��_SV6�EOXCLU-��Xr'ONL�0YY��s<����HI_VՀ�R�PPLYo�RCsHX� �0_M�QПVRFY_I�.Mms$IOv0��}"��1UB���Oj�3�LS����4!���:@�P�$��ĆAUTOCN�E ����.��GCHD�s��_���3sЛAF��CPe�T�!��р� A�o���_�0  �Ԣz�NOCtB$xB�pT��A �����SG�` C� � 
$CUR 8�U��!" �� T@B������ANNUNC�#���䱐b���()%!��-*I&��p@��IC�D @b�`F
"a��POTX� aө�����������[EM��NIߢE��ȷ"�G� A��$DA=Y��LOAD`Ԟ���"��5�� �EF_F_AXI�Fo��%Q�O0<�:�_�RTRQV1G D�a��?0�RK3�0S45 2Fz@]w:1�a�d�A0p/1sAH 0B!�1A�T�2�æ�vDUX��u��C�ABsAIs"�pNSl�1�PID�@PWSsh�5�AWpV`�V_�0|q0�P�DIAGy�sAJ� 1$VX��ET	`�UrT��EJā�{RRf��!�TVE6�� SW|AZ� sP�0�:5q0G}P:13OHP5�1PP|@�SIR|�{RB�P�2�3 %qZQC �BB��H� ^��E`��5q0I��?0����URQDW�EM	SB�?UA�p�EjB�TLIFE�`K#iP��uRN|QFB�U%!zSFBh�a�%"C����N��Y'p�FLA��t& OVڰ�VHE|��BSUPPO(��uRI�_�T��QC_X�d�� gZjWj� g��%!��6�cXZ*�ϡfAY2xhEC��T��DEN�pTBE%!J�� �F_8p��A� @CT�K{ `Q�CACH�*r�bSIZ�V�Pz`�N��UFFI`�oP�ឤ2���62��M;��tL �81 KEYIMAG �TM��!�^q:��Yv�����OCVI9E�@�qM �༠�L~��;�?� 	���р�dNG0��ST��!�r���t����t0�t0�pEMA�ILo����!�5FAUL�"O�r��/����COU��쑁�T���)AP< $d9�p�S�0�0IT��BUF�g;��gE�o�Je��PBe�p�C:�p��:�|�G�SAV�� r�[@�b��@ˇÐ)&AP��p印�D��_e���� �OT겮�3�Pm ��0�z3�AX��#f x Xe�C�_uG|S
^YN_�A.��Q <I0Dk�O�����BM�2�PT�� F!�$�D�I[E7�����R$��$ G���!&�Ǳད�:�9�S�0���-��C_ᰤ�AK�$�����RVq8���DSPnv�PCe�IM��\���<�3@U9��P�] �IP���A�`[�CTH�`3�O�0T��\�HSȓ>�BSC���`e�V��
��#X���*4NV��G;����`Y�e�F|A}�d0>���Z�"�SC%Ba���MER)�FBgCMP)�ET�� TLrFU`D�UY���R�mb�CD R�ܠ'�"���R��
n!UG0*����%��R�%P���C�
ń�-"2��:�o V/H *
�L�� )�9���G ���}�Z {ƥ!{�1{�1{�6q*{�7x�8x�9x�|PTzȄ�1��1��1��U1��1��1��1�ʕ1��2��2�ˑ�2���2��2��2��2���2��2��3��3R��3�˞�3��3��U3��3��3��3��94��61EXT6An!W��߸���V��uş�t���@FDR%D/XTE�V� .�puR�
�uRREM^@9F���BOVM5�*��A3�TROV3�D�T��S�MXb�INp3��PR�"AINDq�BcB
��ɐ}���Ge� �C\�p�UkADO6\��RIVW�R�BGE[AR5�IObEK#�cDN��1`X� zp|`dCZ_MCMp`nuQ �F�PUR���Y ,���?� �P>?o {A?oE� w�1�������Z0*PPM��2@RI��r�ET�UP2_ [ �0q�TDʠ�1p�T�����5�r�BAC��\ T�pr�蔅)�%w#@ó�TIFI�A����d��@/�PT�B�FLUI�t] �@�x;�UR�A���R�Б
���:C_0I�$�S�_?x�J�C9O��"�VRT��� x$SHO^14 #�ASS�-��U̠��BG_ �!.�!���!��!��FORCz#��hDATA)A-^�rFUZ1��]#�2��ˑi�`)A_ �|��NAV=�)�����S��S?$VISI��SC=�SE� ��5UV� O�1&1BFx�4@�&$PO� �I�A�FMR}2��` � ��2���6�!�3J�)�CE#�_����_@IT_Yִ]@�M������DGCL�F�EDGDY�8L�D���5�V���TRH M���sa4�v9? T�FS
��t�b P��RB��}��$EX_RAiHRA1PY�X��RS@3�K5�Fs�G&�	5c �� ֳ�SW��O0VDE�BUG$�A(�GRt� opUz�BKU���O1M� �0P�OZ0Y�@���E�@M��LOOM�9QSMz�0E�� d�����P_E d x�P���TERM[UyedU��ORI֑�`PfdUa0�SM_��`Pg�V�`Q �X�hdU��UP�rig� -���2d��rS�Pe� G�Z @E�LTO���A�FIG�bZ �Agp�T��Tf$UFR��$��aM`ѵ�0OTZgA�TA��lcwNSTאPAT�<�`�bPTHJ�ϰ�E�p�ذbART�؀"e)�؁���REyL�j�SHFTӢ(�a�h_�R��̳J�V �P$�Wph�1p����t�SHI�`�4U � ҁAYLO��m���l� ��a8}!�ޠERV��Sq �x��hgא�b �K��u.�KRC��A�SYM���WJ+g���E��a�y�ұU�א���e@�v��eP��ppE�2vOR2אM3� GRJQ
4jX"�B0V�`G`l�� sHO�6Dk ��aXN� �OCaQ>@$OP�$e��i�����d�ՀRY��aOU��c�PTR�e���|�a�e$PWR��3IM��rR_˃�d0� �P�cUD��c�SV򳠁֔l� �$H�!��ADDR��HMQG�b����ʨ���R�"1m H��S���! ��.�0畞�畫�SEz1�#�PHSܰ
3n $Z À_D��P��.�PRM_�"����HTTP_���H1o (��OcBJ� ��)$���LEyc��d�p � �睱AB_��T@S��S���{�KRLK�HITCOU� À�!퀶������M�SS���v�JQUERY�_FLA!a��B_�WEBSOC�"��HW��a1q�>7�INCPUR�!Ou�ˡ�Č������������IOLN.r 8��R	���$SL2$I�NPUT_PQ$t�ܸP�# ���wSLA�1 sðٿ���s��rNA{IOC�F_AS8Bt$L&��&q�!]�/a�ɳ�@ҳUpHY���lïA�G�UOP5Eu ` X������ā������P������������UQ� M�qqv �l�@;sTAkr��A�TI��.�a�Z0Sն�`PSR�BUZ0ID~0��z���yՏ�!�u�z`w�3��f�G��N��Z0����IRCA��� �x Ĩ��CY�EA{���!���%�R�`�q|�8��DAY_��}�NTVA���i�¦eu��i�SCAepi�CL��������� qy`���ԧb����N_ՀACQ�Ђ�W�rz� O ��������y�G�<]�O! 2y�  ӄ)q{P���P�L�ABzan�Z0t�UN�ISb�PITY0��"ѳ��QIR$6D�|R_URLޏ �$AL10EN��@�� �PH�T�T;_U� �Jt�q} X��t�R��" �0A�D�,J�8FLt@�80�
K�3
�UJR.	5~ ���F|@1w��FgwD��$J�72�O!�$J8B�	7�@\��7s�� 8�	�APHI�@Q��Df@J�7J8�
L_K�E��  �K���LM��  �<��XRK����WATCH_VA�!�pp��FIELDb��y�P&��� �0bpaVyp�ֆCT��E��B`�LG��߁� !��LG_SIZ���@�3@X�O��FD�I� �,Q��]P��� �J&3@J&O�J&�J&�]PJ&�q�E`1_CAM^c�!{@�*h1F���'�$��(�#r��&3@�&O��&��'I�(�(,P�&]P��&�RSI�`  �(/@LN��B�����@{A�g1���K�u1��L~3t2DAU�5EAS�������2�0GH��lQ[�B�OOܑ�� Cr�[�IT8��4<`�n�RE(��8SCRX� ڣs�DIm�SG`nG@RGIPR$D/L@�f�քYB��[�S���Z�W7D[��4f�JG=M�GMNCHH�[�FN�FK�G��I�UF�H2p�HFWDv�HHL�ISTP�J�V�H�P�H�0�HRS"3YHJ��Kc�C4tS �f�x�kG�YUJ��D@jG 3yE�{��BG�I�`PO�WZ&ES�"f�DOC���FEXb�TUI�EI/ ��� /!�dDa�CNc�@��p��� 4	��EpANOGfANA[�ā��AIt瑜��DCASZ���c���bO�hEO�gS?��b�hS�hNHIGN�����A��(��dDE��pTLAL�q��|A��*Є���T�"$���}�h�Ԫ�SA�������ʰ��Z�� �P1
�u2�u3�q���R�`�*І ���V��c ��5�z�x�6��P�6��.�ST��R�0Y���`Q� �$E_�C_�� I�n���8��T)ч Lo��π瀖�x������_�E�NS�_��tD_ �L���X���@���MCh2� =���CLDP��TRQLI��D�2�FLGZ�2�3�f�b��Duf�`�LDf�P�f�ORGjQy�~�(RESERV���Ŕ��Ŕ� #�3�� � 	O�jUA�Ff�SVX0D�R	����'�RCLMC�5�şןG���'�pM�ՠJ�/�3$DEBUGMAS�ÐS�D�"��T�`p�E�� TZ�
�MFR�Q��� � ~�HRS_RU���ځ�A)��UFR3EQ� J�$``�OVERh����v�|P�AEFI���%������ӡ�� \ ��$U���?����P)S�p7 	�C�06��BҒ�G�U�Н�?�( 	"MISC�i� dq1�RQ�5		TBB@�� 1��aa�AX9�!|	�"�EXCES��c۳M��.����9���ܲSC� O� H���_G�@��,��� �2��K��a�|��B@��B_��FLIC��B@QoUIRExSMO��yO��d��ML܀M��� 
��19����5�`pMND�1e�/�o2f2�x��D�#�4INAUT(A�4RSM� ��p�NZ�b!�S^�`0e�PwSTL.� 4��7LOC�RI1P�;EX��ANG�b��n��ODAե��1p�x MF�% 7�+�ۂ|@�e�c0��gSUPᅠqFX/ �IGG�1 � ���ۃb!Cۃ�Vۄ ��V�P���R���R���`���SD�w��TIjȯ��b!M ��� Mt-�MD*��)8��`C�L�@�H�C�GDIA�D�2 W]APC��q��C�D�3)3�qOh�/� a�CU�V����"��OPA_��.� �`t �7㉠f��
 B��P��>P���P���KE�RR�#-$B8�����ND2N�N�D2_TX�XT�RA�cp`��9�L�O�0/�_��	�i2����k��RR2൜� �-��1A$� d�$CALI��c%Gt�a�2�pRIN�!��<$R� SW0�S� `�ABC>�D�_JV ��� 7�_Ju3K
E1SP�$��� PEl3k����� �J`��撚�OiqIM`�ŲCSKPS��� �c�	J�1ŲQ�%�%'�_AZ#��=!�ELNq�N�OCMaP�Ʊ��z0RT���h#�1����1ћ�(o`�*Z�$SM�GMP�n�JG�S�CLB���SPH_@�`Ű+0�#\ � � ORTER��`R� _�`�*�AP@�G�Ų4DIS!�"2[3U�DF�p<1�LWB8VELD�IqN�Z`e0_BL�`��m4���J]4r7�7��4�pIN� �������5QB��
�1��_̰ ��5�2#5l���4z�936ٰDH�B�r ����p$V0� ���#oa$� �l���$\���ൡH �$B�ELN ��!_ACCEs1 �H`��@OIRC_06����NT��/�$PSB�7�L�p��DL� �0�G3�`�F;�I�GD�C�G3�B��E�_�q�PB-P3Q����A_M�G��DDPQ2��FW����ClU�C�BaX�DE�[PPABN6�GRO� EECR�q �_D�!�q�����A�p?$USE_� �c]P�CTR�dY�P�b@"� ��YN߰A a`f�Z�aM����ĵbJPO_0�AGdINC���RpT�ig�.�ENC0L񦲰�A�B��@IN7�I0�B�e��$NT]3�5NT23_@2���cCLOQ0���`-�IP� ���fF0����� ���e��C�0�fMOSI�UQ����3Q�ŲPERCH  s+�2 ]w�hs��rn���@c'["e
P2P�A�B�uL�T�����e��8z�vvTRK�%ʁAY��s��,��r;��0��n&��wbȠMOM��»������S��G��C�R� DU��(RS_BCKLSH_C�r����<v ,�"c��݃�b�1a%CLALM�d��m�@�CHK��NGLRTY��5�d�����_Z�1t_U	M��l�C��^Q�!��n��LMTh_L��V#��j�E��Ð�� ���E���H}���r�&�xPCnq�xH���TUl�CMCv^PbWCN_�Nuc��SFtA�yVb�g��!8��r��<�CATs�SHZ��bT�f]�����f��A�	� QPP�As�gb_Pr�V�_ �� 3�Qp�C�U�F��JG>�X�I�K0OG|V�2TORQU�P �/sL��P��Gr1�P��_W��,��!QAٴPBCصHCصI�I�IHCF$�˱�-��ZPVC�@0����N��1T�RPh�$!Z�JRaKT̙ƴ�DB� �M���M��_DLBA�rGRVߴ��BC��HC��H_����@��COS�p �LN��6�W�=�B@8ٵ @8�
�t�b�(���Z1�Gv��MY?Ѳ��=|'���THET0uNK23HC��<C@�[CB�CB<CC� AS�'�
�5�BC5���SBBCS��GT	S��QCo/��'�x�'��q�$DUC�@�w���t5��5Q�qY_��NE��AAKS�z)!8 @��A����'����LPH����e��SW�o�b� o�q���֙�����EV@�V5�2@X�Vg�UVt�V��V��V��V��V��H@�Y�_PW�ܡvt�H��H��UH��H��H��O1��O@�O�	V�Og�O�t�O��O��O��O
��O��F��"�~b���3�SPBALA�NCE_�ѮLE6j�H_��SP�1S���b��q�PFUL�C�"�"q��:1=�|!UTO_>�F��T1T2B)�B2N %��B�`b$�!f� ��(�B}C��T�pO50�A>ɰINSEG�B q�REV�& p�aDI�F��91��'321�	�OB�!	��Ó��2���`0���LCHgWAR�R7BAB%�~��$MECH+���9a?1T�AX9�P��X6�#B7 � 
pY2��{A�eROBQp�CR�r�5M� ��CyA_A�T �� x $WEgIGH6`�$1�d�3X�I6a�`IF�QNjPLAG'b�S'bܲ 'bBILEOD�o�#p�2ST�@�2P�!	��0`@Ơ�1�0���0
�`yB(aA� � 2�.t�6DEB�U�3L�@<B��M'MY9�E� N��D��$D�Axq$��@S���  ��DO_�@A�1� <�0VFL U�(a�IB&B@N�c�H_p�(`�CBO� �/� %��T�`�a⊑T�!~D�@TICYK�30T1�@%NS���WPNQp1 �CQpR�Ԁ(a!2iU!2uU�@P�ROMP6cE� $IR��&aL�8�R�p�RMAI��aa48b�U_@�S� tB�:`R��COD[CsFU.`�6ID_pp�e� �R�G_SU;FF
� Ca�QdRDOlW� mU @lVGRC!2Id�S Ud!2`e!2le��Id�D�e@��0H� _FIvZA9�cORD&A3 �0�B36��b|&a�@$ZDTe� 	
CA�E�4{ *�!L_NAQ�WPriUDEF_I )xr�V5tuU-BhV7D`hVasuUou�VIS��@���A��hT�suS3tD���D4l���7BD5 (���t[CD��O��BLOCKE�Cci_`{_�W�qIbC`UMHe rIdasIdouId�rUb K�TeDsUdtUb5F�� �q`c,0B�`er`eas `c���EhPP� �t,P�q��@W*�)� �	 �TE���D� ALOOMB_C�^�0�2wVIS!�ITY�2�AS�O'CA_FR1I2#��� SI�q��B�RTP��_P��3tC
�2W��W��������9_��jaEAS�3jb@d������p�R��4���5��6�3ORMU�LA_I��G�	w� h �N7��ECOEFF_O ;Q� ��;Qr�G��3S�0�BCA �O�C�CAGR�� � �� $ �u"�BX+PTM�� �AR(�,%��CER� T	�tn�`�  +"LLkd:�pS�_SV�tw�$L��`���v��`�� ��SETU�sMEA�P(`F��0�CA�b�0� � ���0 �@o��Q2��q�rWP�q�	�tբܑubÕQ��p�q�p+���� ��PREC�a� ? �MSK_���� P�11_USER^!�"}�0��}�^!VEL"�}�0ȥ�!1I�`J �M�TQCFGs�� � YP� OG2NGORE�0P���0~��� 4 ݳ8B7�2H1XYZ�cJ!�o yC�1��_ERR��1� �I�Q�P�ۣ@�aAi����@B�UFINDX� �;�MOR� H�0CU@�QH1����Q�a���"�a�${0��~q����;���G� � $SIj����P��!��VO����0O�BJE���ADJ1U�B�� �AY�p5��D.�OU�`Վ�\'a�b=��T� p]��\��BDIRa��i�� ��"�0DYNH쒣2��T6 �R���,P&@��OPWO}R�� �,�@�SYSBU �SCOP��cҎ���U��b� P ����PA�����C2�OP^`U��!��!XB�AI�IMAGS��0U�7B3IM��o�IN��@�~n�RGOVRD��	��K�PM�m�0� P߀�s��H2L�B=�|� �PMC_E�`cъANM��A�B11�B�@��SL�t��� ��0OVSL:�&S�DEX�q}p"/2G2� ��_��G �`��G�`Qfa�B�C�0p�%�c��/_ZER�����s�� @вb5O&`RI��s0
��P��	��qPL�Ĵ�  $FRE�E��E�������!�Ls����T<D0;@ATUS㰤AGC_T��r�UB� _H��s�A4�`t��� D�AI�2RL���a2S�an S���X�EY������ �0XUP��p�qCPX�PF�D3��^� �PG�Ÿ��$SUBGb5���G�JMPWAIqT�V_%LOW�8BQ��@CVF�QZP�G2b!Rz���U3CC� R��MR�'IGN�R_PL�DBTeB;@P�qH1BW�Pd�$��UP�%IG0�z�PIG3TNLN�&"2R�����N�P)�PEED�8HA�DOW;@�����E�7S4F1!4pSPD.s�� L�0AV�5ps0�3UN�0"+02!R��LY�`� �Q���P��v1��G�$��M�P�@L\+�NPA�T�2�xD��PIP%w0�>��ARSIZ�T���c|q�Om`�h�A�TT���"\�B$�M�EM�B�A>C�3UX���e�PL`�ļ� $���SWIT�CHZ"�AW��ASr�B�BLLBv1��� $BArZ�D�s�BAM� h���I��@J50�����B6�F�A_KN�OW�3R��U!�A�D�H۠~0D��5YPAYLOA鱱�SS�_s�\W��\WZYSL�A�mpLCL_�� !���R�A����T���VF�YC�K��Z貓T��I�XR�M��W_ҬTB���JL)a_J�Q����AND^�9�8d�R�Q����PL�@AL_ ��@~0���A��k�C"�DXSE!��sJ3M`af� T���PDCK��r�C}OŰ_ALPHqc��cBE��W�qo�l ��Т�!�� � ��40R_D_1YZ2�TDŰAR�4x!uxEv0s��TIA4_yu5_y6"�MOM��@ks�sxs�s�s��Bv �ADks�vxs�v�sPUB��R�t�uxs�u��r�Fp��� L$PI�1s��^WP.��xY.�I:�IH�IV�<p}Q7��!�� !��b�ӆ��73HIG�C73w%p4І p4w%� z�І�߈�!x!w%SAMP����B�ЇC�w%�@>c 5�q���7 �Ҁ�  ��p0"p��0p�������hp���	���IN ќ�&�ؘ��ϔw"ښ����:�GAMM�ƕS[%�$GE�T��o��D�d��
�ϡIB��2I0�$HI�_��sЩү��E�м�A��٠ʦLW�����٩�ʦ�b贆0caC�%CHKh��� 	��nI_%� ����\bxΑ�����s����v���c ��$�h 1���I>� RCH_D��'� �$)�LE��������hذ�0MSW�FL�$M�`SCRF
(75_����3�� dƧ���kp��x�p0�����SVv1�P���v�Kǿ�	���S_�SA�A�����NO�`C���d���� d_v_\�J�:ۂ�+R��w�0sD<�4���40�� zʴ�ʈ��چ�1��� �ՕәS�Ak0L���� � ��YL,�a������-��� -���b��9�az�HK����W�{����py�Ȳ�M� ��P��`a�$ 7��"r�M���� � �$���$W���ANG]�Q���d���d@���d��d� נNPP���C��ϐX�0O�c�ΑZq��� �� -�<�OM��"���1�C�U�g�bpCON���0}C�a_�B� |�a�����y7xs7 �s��dzdO~z�A��� J���Ǡ �PP A�PMO�N_QUG� �{ 8�0QCOU��nǀQTH� HO&�n� HYSD@ES�BF� UE� ��@O5$�  �@P�৥���RUNZY�0 O��� � POP+�%����2ROGRA(��x@:�2�Ov+�IT�xINFO��� �A_��8�ȫ�OI�� =(ʰSLEQ�����b�S_ED�d � � ���r�KԙQI#��EȠNU�'(AUT��%COPY�Q��8,����M��NB F+U�PRkUT� I"NF2U�B$G0�$Xa�PRGADJ!�fBX_��2$�0(�&~��&W�(P�(���&73� �NH`_C�YC���RGN�SD���LG�Ob��`NYQ_FREQ�rW����^1RD)L�P:BV0�!�s���CRE���c��IFH�jNAK��%�4_G�STA�TU å�MAI�LI�S&@V��ǀL�AST�1�a04EL�EM:1� �EaN�AB�0EASI &A��v�n�?�B���GF�����I���U2`���� �|BAB�C	PRS�LV	A�Fa��I���qU����JP�'c�FRMS_TRvCΑ��Ci�����A�D E���& 	SB 2�  �V��9V(b8WR���RNTdW&�
�DO`�P�W}�
�22PR �z;0��GRID}��BARS��TY�'C��O�p!� _�4!� �R�T�Oo�74� � |� PORXc�.	bSRV�0)(d fDI��T!pAaTd���^g��^g4\i[�^g6J\i7\i8@aFj��:1�$VALAU�C��9D��F65�� !"E��lb�S�1��_@AN����b�1R c17ATO�TALH��qCsPW�K3I�QYtREGENWzlr�X�H@c5v� TR�C�WqC_S���wlp\CV�!p���u���1GRE�3��P�6B+.  sV_�H�PDA���p�S�_Y�i�o6SV�A�R��2� �"IG_SE�3�p b�5�_/�tC_�V$C�MP���DE�M���Ie�Z��^��zF�HANC�O� p&Q$E�2���INT?`iq��yF%�MASK=�.�@OVR�P� �P ��1Α�W!��T� 4� �_XF�{�V��PSLGV�:1� @K��p5a���Ap�JpSh��4��U0>�!����TEa��`G���`�U�Jd�<��3IL_M~4���p� TQ� �����@-�\�V4�CB�Ph{�4AL�Mc�V1b��V1p�2�2p�3*�3p�4�4p�����p:����p��j�|�IN�VIB��<�)�T��0�2,�28�3,�38�4,�48� hR�ґ��� �T �$MC_F�  ����L����ׅ7pMb8�I׃���S ( ���n�KEEP__HNADD��!�$�@��C��0��Q��?��O��| ��p�p�܇�REM'�IqbL�c�h�U��4e�HPWD w �SBM�~�PCOLLAB���p��5q�2�IT�50`�w"NO��FC�AL��� ,��FL�A$SSYN���M� Cq���XpUP_DLYz!�DELA?дJq�2Y� AD����QQSKIP��� �`-O;�NT�]�i�P_-V�� ^U�*����q���q�� u`�ڂ`�ڏ`�ڜ`��Щ`�ڶ`��9�!�J�2R0� �L�EX�@TX3N�7AN� ��N�}� RDC���� ���Rz�T#OR� ���R�1��x���;TRGEA�r8h@��RFLG�^��5�ER���SPC��1UM_N��2/TH2N�Q�A�� 1� ��A��Q62 � D�Kш��@2_PC�3]�S���1_0L10_C}2��2���7 �� $b�  ���	ViR����0�� �\Ub����m8rj��C1��*=��ID� Gy�XUVL1a�1n��� ;10c�_DS�����<��P�11!� �l�����#C��ATE��$�Q���f���;T�3�HO�ME�� f2n�t������3n��'9K,0f4n�n������ f5n���/!/3/E/
�6n�h/z/�/�/(�/�/�7n��/�/@	??-???c�f8n��b?t?�?�?�?�? �fS���!�  �Ag�p��;�zc�Ed� TC�tD:vtCIOꑔIIt@f�O��_OP�E�C4rlC��POWE�� ^@�l�q�`5�5s ����B$DSB��GNA��3s:�C��b0��S232zE� ����5���ICE;US=sSPE(��a�PARIT �2qO�PB���bFLOWFO�TR9@?rt�UX��CUuP���aUXT���a�ERFAC�ZTT�U.p �2PCHa� t�఩�_`Py���$L ��pOM8���A��8�𥀯�UPDư��f�qPTU@��EX��8#hc�EFA8�����BSP�P�a��|�`�7$USA�X��9��EX�PI��$(`�pY�eR_$�q�`mQ�fWR�OI�D���f��FFRI�END��L�$U�FRAMc�pTO;OLvMYH��r�LENGTH_V�TE�dI�;s��$Z pJxUFIN�V_^ ��_ARGuI%���ITI��bBwX�Sw�vG2�gG1�aꀎc�r�w�_r�O_XP��L�+q4���N�Sc��Cp�Pr�q��G���Rǁ󐒧�XQ؂��h�U���U�������PUd�X nm`E_MG`CT�c�H��h���U�dScG��W�`ć��لD]и@KȅJӂй�������$-� 2!���an �i1�h�`U2�k2=�3�k3�j -����iK���F�`l�P�`x�|�NtV�uV�ТPqC,��r�P��� �V������R��pr�.���E9�<�Os�)E$A��T�P!Rh�U�k�ǓS��P����Sb;Q� ! �ႃ"��K��"����S`�p�p��
 ��$$C��S�������9�9� }ؠVERSI�`����i���I#PP��AA�VM_�a2 �� 0  �5�V�b��S��� ��	 ������9� �����ζ����ϧ��0R�d�l�0�BS^ r�1�� <@ϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� ����������'�9� K�]�o����������� ������#5GY�k}����|�C]C`XLM�@�����  d�IaN����qEX?��2_`=� �9��0�IOCipq ��PZXQ��{�IO'PV 1]=�P $-��ұ0�!̺ �?���  ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{���ϟϱ���� LAR�MRECOV �I��LMD/G �����_IF  ���p߂ߔߦߴ��^���������, 
 �G���� m�����$_��� ����� �2�D�V�h���NGTOL  �I 	 A �  ����� PPI�NFO %�� $������  1�I
�8r \������� &W�p�Rdv �������/�/*/x�PPLIC�ATION ?�����LR Han�dlingToo�l y" 
V9.10P/25���5'
88340�z#�*F0�!�/13�1y#�,�/�"7D�F1� 5,y#Non}e5+FRA5/� 6�-B&_A�CTIVE��  �[#��  X3UT/OMODb0)���U5CHGAPON�L�? �3OUP�LED 1M��� �0�?�?�?O;CUREQ 1	M�W  TILL�	XOiE_ ~D�;B�m%MD�H6E�2cJHTOTHKYwO��D\COUO_�O7O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_oo#o 5oGoYoko}o�o�o�o �o�o�o1C Ugy����� ��	��-�?�Q�c� u�����󏽏Ϗ��� ��)�;�M�_�q��� ���˟ݟ���� %�7�I�[�m����� ��ǯٯ�����!�3� E�W�i�{���翱�ÿ տ�����/�A�S� e�wω��ϭϿ����� ����+�=�O�a�s� ���ߩ߻����������'�9�K�CETO��d?X2DO_C�LEAN�?V4��N�M  �� �O*�<�N�`�r�ND?SPDRYR��U5HI�0�@����� &8J\n�p���R8MAXI  ��|�~A�7�X���!��2�!X2PLUGGp�0���3t5PRC��B�����.�O3����SEGF�0Kz�������//&/^�LAP����Cz/�/�/�/ �/�/�/�/
??.?@?|R?�3TOTAL�|�3USENU���; ��?~B@R�GDISPMMCʚ�AC��@@$���4O�����3�_STRING �1
�;
��M�0ST:
)A_�ITEM13F  nT=OOaOsO�O�O�O �O�O�O�O__'_9_�K_]_o_�_�_�_�I/O SIGN�AL-ETry�out Mode�4EInp�PSimulated8A�Out�\O�VERR�� = �1007BIn �cycl�U8AP�rog Abor�c8A�TStat�us6C	Hear�tbeat2GM?H Faulug~cAler�i�_�o�o �o�o�o $6H ��/K��AOK �������� )�;�M�_�q�������p��ˏݏ_WOR� /K���=�O�a�s� ��������͟ߟ�� �'�9�K�]�o�����PO-Kia��-��� ܯ� ��$�6�H�Z� l�~�������ƿؿ����� �2ϴ�DEV ��]�ЯJτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶�����PALTu}�-� ��)�;�M�_�q��� �����������%��7�I�[�m���GRI � /K���������� '9K]o� ����������0Ru}I��#q �������/ /%/7/I/[/m//�/x�/�/7PREG� � a�/?'?9?K?]? o?�?�?�?�?�?�?�?��?O#O5OGOYO�]��$ARG_�D �?	����A��  w	$�V	[�H�]�G��W�I�@SB�N_CONFIG(�P�K�Q�RQ�A�CII_SAVE�  �TQS�@T�CELLSETU�P �J%  ?OME_IO�]�\%MOV_HVPi_o_REPL�_�JUTOBACKAQ��IQFRwA:\�+ �_,�&P'`T`�'h�� k
P �18/02/�09 11:06:04�&�H�-{o0�o�o�o�\���o@%7I[�&��o ������n� �+�=�O�a�s���� ����͏ߏ�|��'��9�K�]�o���X� � �Q_�S_\AT�BCKCTL.TM����ҟ�����[INI�AeV�S?MESSAG!P/��Q�@SQD�ODE�_D[P$VUb�Ox_�q��SPAUS͠� !��K ,,		��@�Eѯߧ ů������Y�C� }�g�y�����׿��ӿ��������TSK�  ��o��PUgPDTh�-�d~��~�XWZD_ENqB-��J��STA,���A~ŎAXIS�@U�NT 2�EQ�P� 	D��p���� &~��X���?H�F�*�� ��  	X$U/k�>��-~�  ��U�X;`UX�T����Pߊ�����METrK24�-S P���A�AK]*�A�{/6�1�Ad�
A;L���75n�8��S8cff4�D�D7��6���@��SCRDCFoG 1�E�Q' �)UR�߆�������o�*Q %Ys�0�B�T�f�x��� ����������`,�����G�QGR���r���k��NA�P�K	�Th_ED�+�1V�� 
 ��%-��EDTA-Y�Z�M�
T�zP-�S��*�B��otV��  ��u2~�[\���'��/Yk/�w3 J/��/��s/�/%/7/�/[/w4?�/c? �/�??�?�/?�?'?w5�?R?/Ov?�O@vO�?�?eO�?w6�O O�OBO��OB_�O�O1_�Ow7z_�O�__ ��_oU_g_�_�_w!8Fo��o��oo@�o!o3o�oWow9�o_�o��;��o0�o�#wCR}�_ *�<��]�p���_���k � NO_DE��yk GE_UN�USEu�IGALLOW 1�	�   (*SYSTEM*���	$SERV_�GR��*���REG�3�$U���*�NU�MX�}�k�PMU>�LAY�С��PMPAL|,���CYC10���ʞ�����ULS�wѭ�G�̒��5�L��?�BOXORI�\�CUR_,�k��PMCNV���,�10����T4D�LI��%�G�	*P�ROGRA2�PG_MI������AL¥����B��*�$FLUI_RESUЗX�b�
����������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯�������H�k �LAL_OUT ��T�WD_ABORѐ��jO��ITR_RTN � st��O�NO�NSTO� z� �b�CE_RIA_�I��z�������FCFG �
��s}��_PA�9�GP 1����Q>�P�b��!�C/�����z�C��C ��(����C�8��@��H�� CUX��`��h��p��Ux}�������������	su�?���HE��ON�FI��Y�3G_P6r�1�� ��ă �}������|�3KPAUSI�31`�� ��� C`1oU�� �����/5//�Y/k/Q/�/Mo�N�FO 1`}�� � 	-���//�� �"�DA��/?������µ�B�QK��� D��b����B���B�3�0S��B��� 0²��B���j�r�7�5B�ai�80��O�����swV2LLECT_����&A���~7E�N z���2W1ND-E�3�7eヂ�1234567890�7~rD����?��6ss
 ���q) 9O^OD�8OJO�OE�|O �O�O�O�O�O/_�O_ _w_B_T_f_�_�_�_ �_o�_�_�_Ooo,o >o�oboto�o�o�o�6vB�2�; �=>�2IO  �9�1�yxy�as��/wTMR�2!}�� Jy1
�o�~> ">}�z����9_MORr#
� �'	X��!X�p� ^���������1� �q�$?�,C?,,���/�K�TqJr��P[2&�?"�+�a�s�����
R���t7���u��y���5���ss ���9PDB/��(7��dcpmi�dbg�]�v o�:���nD�pI���m�/  ��nG�毆���ï��.�����mg�x�C�Ů�fg����-ſ�`u�d1:���z'�D�EF 'y(Is)���c�buf.�txt�g��%�_KMC8�)7�!sd����7�*��������|ƟCz  B3A� C�lCyC�d;�p������-D���D���D�J0?M��D�I�D���~�-F���F���F�U�CwH�S�F��P*����,|��t7A�pH �pJH �H ��t
����� E�@ Da � D�  E	�� D�@ ��;��| Fp F"�� G=�fF���G'i�-G�>�Gg� G�K  H�<=H�&HyMc���  >�33 ' `C/��n)��F�5YT娂��A��|�=L��<#�� �Vq����ξ��RS�MOFST %x8ʝ/P_T1���DE -3�����q��Tq;�������?���<��;��EST2�+8�PR�2.a?����+C4���|���p���������C��B�f��C����H���p:d� ���T_~2�PROG ����%x�V$INU?SER  �5(�$KEY_TBL�  �"�	
��� !"#�$%&'()*+�,-./�7:;<=>?@ABC2��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������0�������������������������������������������������������������q* L�CKt��&t ST�AT���_AUT/O_DO�6���GIND�4�V1R����T27/�STqO@/� TRL, �LETE�7~*_�SCREEN �?�kcsc��2Uo MMENU� 1/.� < ED?[�/?J?ճ '?M?�?]?o?�?�?�? �?�?�?O:OO#OpO GOYO�O}O�O�O�O�O �O$_�O_Z_1_C_i_ �_y_�_�_�_�_o�_ �_oVo-o?o�ocouo �o�o�o�o
�o�o@ )vM_��� ����*���9� r�I�[������ޏ�� Ǐ�&����\�3�E� ��i�{���ڟ��ß��Ϲ�#_MANUAyLs/�!DBCO �RIG�'�/�_E7RRL2 0��a�aN�����ǯ P��NUMLI;�Z!�����
P�PXWO_RK 11�����'�9�K�]�o��DBwTB_�! 2���ç����DB__AWAYX�a�/GCP ��=E�ö�_AL;��òT�Y�r �%��I�_r� 1}3#� , 
�`T��B�ω�_M �I��Ѽ@����ON�TIM�'���ɼ���
�$�MO�TNEN��z$�R�ECORD 19Ξ� ��ψ�G�O�O�=߈�Ҳ{ߍ� �߱�Hع���O��s� (�:�L����߂��ߦ� ������� ���$��� H���l�~�������� 5���Y� 2D�� h��������� U
y�Rdv ����?�/ /*/�N/9/G/�/� �/�/�/;/�/�/q/&? �/J?\?n??}?�?? �?7?�?�?O�?�?FO �?jO�?�O�O�O�O_O �OWO_{O0_B_T_f_��OòTOLERE�NCдB��ްL���P�CSS_C�NSTCY 2:J����i_���_ �_�_oo'o9oKoao oo�o�o�o�o�o�o�o��o#�TDEVI�CE 2;�[ ��vu���������*��ϭSHNDGD <�[��Cz|{�TLS 2=]}<�����Џ�����>��RPA?RAM >0� ���|��}�SLAVE� ?]�I�_CF�G @J�*�d�MC:\�PL%04d.CSV)�b��cџ�RA ��CH�o�o�*��F��w�*�6�c�s�xa�`��JPѓ��|����r�_CR�C_OUT A�]}��.�_NOCO�D~�B0���SG�N C&��&j���21-A�PR-21 00�:38�*�0�9-FEB-18? 11:06��v LIX�v��r�*�s�Iu5��M��Þ��������VERSION -��V4.2.1�0��EFLOGI�C 1D�[ 	��+�ɘ�!���PROG_ENB��e�A�ULS�� �d��_ACCL{IM���������WRSTJNaT���*��MOJ������INIT cE�Z&�*� ��wOPTy� ?	�����
 	R5�75*�+�740�6J1�71�5�[�1U��21ԋ����TO�  ݉����V.��DEX��d��p����PATH ۦ��A\��9�K���[HCP_CLN�TID ?Ѷ��� ��"S��QI�AG_GRP 2�J�� Q� 	 @K��@G�?����?l��>��������Q �������P)��?�b�?�PT�i�^?�V�m?Sݘ���f403 6789012345{������� ��s���@nȴ@i��#@d�/@_��w@Z~�@U/�@O�@I��@D(���𷡋@���p����PAe�P�P�B4��jp��ط�
��1���-@)hs�@$��@ bN�@��@�����@�D@+����������	 ���R��@N�@I�@D��@>�y@9���@4� .v�@(��@"�\P�bt��L��@Gl�@BJ�@<z�@6��0��`@*� $N?�@���� $=q@����F@|��@33@��R@-?����?��`?�+hz����Y"�J�-@&��@N���!�?�?� � �//*/</�-�/ ?�/&?8?�/?Z?�? ^?�?�?@?R?�?�?O �?4OFO�?VO����@9�Q�i @��V���AY����?��z��A��5AF��A4��@��L4�R��A��@�p]� R�Q�R-P�P��@�� ��Ah���=H�9=Ƨ�=�^5=�>P��>���o=�,d_�,P�� ���C��<(;�U\� 4���ඨ_����A@��? ��pO�_xM�_o0o�� �T<ofo ovo�o~o�o��o|I>��y�b��R=���=���zq���G�G��� � ��!�!��NUt@�T��V���uB�� B��B��B%C�����~'����u���q�q6|䏁\�&���g���)PB�3pB�B A�@��"���m���<~��  3��T��40�T�����g9y�fw�ڔ�����D��\��3aB��Fp�l���r�ݏȏ���x�"�������3�����B?���?�Ǐp� 돔������ܟ�9Q��0T<��I;�����������XѶ�E�=����CT_CONFI�G K�m��eg7Ų�STB_F_TTS��
Yɠ��Ȱ��������M�AU��N�N�MSW�_CF\�L��  ���OCVIEWf��M��ᄀ�� A�S�e�w�������/� Ŀֿ����ϭ�B� T�f�xϊϜ�+����� ������,߻�P�b� t߆ߘߪ�9������� ��(��L�^�p�� ����G����� �� $�6���Z�l�~�����,��D�RC�N(E��!P�����!E4�iX���SBL_�FAULT O�����GPMSK����P�TDIAG� P`��qo���o�UD1:� 6789012345t�n���P*�Sew��� ����//+/=/�O/a/s/2���R
�B�/J�TRECP�
?)�+A >?P?b?t?�?�?�?�? �?�?�?OO(O:OLO�^O�/�/�/�O�UM�P_OPTION����ATR袒��	��EPME���OY�_TEMP  _È�3B�5P9��TUNI͠���5QܦYN_BRK� Q��EDI�TOR�A�A_�R_~� ENT 1R���  ,&M�AIN��-�OdM&�PICK�_o &DROP�_�3o�PPROG_�#o`o&}�os��to�o�o�o�o�o �o/SeL�p ������� � =�$�a�H�p���~������ߏ�؏����PMGDI_STAHU�$�5Q}UNC;�1S� �dO��v��N
�Nd�Oݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W��En��������� ʑ��ؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@ߺ� g�q߃ߕߧ������� ����%�7�I�[�m� ������������ �!�3�E�_�i�{��� ������������ /ASew��� ����+= W�Es������ ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?Oak?}? �?E?��?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ G?Y?c_u_�_�_�?�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7Q_[m ��_����� �!�3�E�W�i�{��� ����ÏՏ����� /�IS�e�w������ ��џ�����+�=� O�a�s���������ͯ ߯���'�A�3�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �9�K�U�g�yߋߥ� ����������	��-� ?�Q�c�u����� ����������C�M� _�q����ߧ������� ��%7I[m ������� !;�EWi{�� ������// //A/S/e/w/�/�/�/ �/�/�/�/??3!? O?a?s?��?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_+?=?G_Y_k_!_ �?�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	#_5_ ?Qcu�_��� �����)�;�M� _�q���������ˏݏ ���-7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����%� /�A�S�e��q����� ��ѿ�����+�=� O�a�sυϗϩϻ��� �������9�K�]� w����ߥ߷������� ���#�5�G�Y�k�}� ������������� '�1�C�U�g��ߋ��� ����������	- ?Qcu���� ���m��);M _y������� �//%/7/I/[/m/ /�/�/�/�/�/�/�/ !?3?E?W?q{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O?�O+_=_ O_i?__�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o __#5G�os_} �������� �1�C�U�g�y����� ����ӏ��o�-� ?�Q�ku��������� ϟ����)�;�M� _�q���������˯ݯ �	��%�7�I�c�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ���������� /�A�[�M�w߉ߛ߭� ����������+�=� O�a�s������� �������'�9�S�e� o��������������� ��#5GYk} �������� 1C]�gy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/I�??)?;?U _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�/�O _!_3_M?W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�O�o+E_ ;as����� ����'�9�K�]��o���������ɏ�o ��$ENETMO�DE 1TFu�  �`��`�e�"��R�ROR_PROG %��%�fe�r��@�TABLE  ��P��ß՟��@�SEV_NUM� �  ��	��@�_AUT�O_ENB  �,��=�_NO� �U��!�� W *�]��]��]�	�]��+\�v������6�FLTR"�4�H�IS��a�/�_A�LM 1V�� e��d]��`+���6�H�Z�l�~�����_\��<�  ��[��"�պ�TCP_V_ER !��!]����$EXTLOGo_REQ֦�-��'�SIZ0�"�ST�KM�K��$�T�OL  �aDz�ޢ�A "�_BWD��������'��ûDI�� WFu��� ��a��ST�EP�������OP�_DOo���FDR_GRP 1X����d 	пm�"�^��n&���c�?��$,�MT� ��$ �����^ӳ����^�B��%BZ���B�S�B�ȟ�B=�����(UB $B��V�Ae~�A�?�A������� :�%�^�I��m����  AJAs?�Y>(�����`
 E�� 	�<���a?�{��������?�*�c���A@�����@�33@�������@���L�x����^�F@ ������������L�F�Z!D�`�D��� BT��@7�����?���O���6���u���5�Zf5�E�S������J�ƿ� .H� ���X[x��n4�x�FEATURE� YFu��&��LR Han�dlingToo�l ��bEn�glish Di�ctionary��4D St� a�rd��Anal?og I/O#,�gle Shif�t?uto So�ftware U�pdatedma�tic Back�up�	�ground Edit� ~�Camera:�F>Common� calib U�I��n��Mo�nitor�tr~� ReliabS��DHCP��
D�ata Acqu�is�%)iagn�os�7?+ocu�ment Vie�we"''ual �Check Sa�fety��ha�nced��
�%s� Fr��xt.� DIO �fi�u$�'end� ErEr Lt"	=�'s9�r5�  ���
FCTN Menu� �v##[7TP In�J0facq5�Gi�gE�>�5�p Mask Exc� �g�'HT�0Pro�xy Sv�$�6i�gh-Spe� S�ki��6m � mm�unic�onsHurh0J0:/;�2�connect �2:Hncr�0st#ru8Ja@e�!� �Jt%�KAREL Cmd. L�0�ua�8�CRun-;Ti� Env�HK0�el +�s�S�/W�Licen�se�#�,0Boo�k(System�)�
MACROs�,�2/Offse�ZUH� w8/"PMR �s.M}M@!�l�,MechSt�op�1tQ@Y"Ui2V�Vx� 7�L^�odTwitch��_aSh!.BV�[OpctmoaS�0fi�^�aVg0GUulti�-T�0��	PCMO funkG�ia�P�tiz~h�goV$R�egiPr@�fr�i� F�k�f8Num Sel�U�i�  Adju@�n q<V1}tatu�aI��*�RDM Ro�botscov�e�ueav`� F�req AnlyNGRem�P�!n|�u�rServo� ��P�SNPX b��B[SN�0Clix�!�WLibrD(��  �T:��vo�@=th0ssag~e��� l5Q&�/I|�=��MILIB��~��P Firmu:��Ph3Acc���TPTX4/��el�n5PǏ���1U��o�rquTimul�a!�E�u�PPa��A���!!c&�0e3v.��mri� ��USR EVN�Tğ֐nexcept� �pn�#ѕ�(@VC�rBB�X�VU 6��G�:�A�S��SC�y�SGE쎯��UI&Web Pl`vǮ�q0O���0�$�!?6ZDT �ApplD�
iP�0a!�:� Gri=d�qplay=����W�R-�.��h!�N��B^P}200i<V4+scii�1r�Load� �Up�l���f@I�Pat�V�ycS�B�`��� \6RL��� ۩�5�MI Dev�@ �(�qR�f�?�gss�wo!�_64M?B DRAMM����FRO�Ͼell�:�sh��#�c�.k �rp��5�tyBSs
r7̬r'`.?+`�p�!"=-o� 2�=a5port�.�p4�r q�-T1 �{x]P��No m�p�c$筴OL��S�up��Fa�hOPCg-UA�l�T �2�eϓ�S0�0cro�a|�s:����~���uWest�uS��e2'texV��up�1�#Ɣ�PP�00�oVi�rt�!�sR�std�pnÛ�� SWI�MEST f F	0����������� ������ MD Vpz����� �
I@Rl v������/ //E/</N/h/r/�/ �/�/�/�/�/??? A?8?J?d?n?�?�?�? �?�?�?O�?O=O4O FO`OjO�O�O�O�O�O �O_�O_9_0_B_\_ f_�_�_�_�_�_�_�_ �_o5o,o>oXobo�o �o�o�o�o�o�o�o 1(:T^��� ����� �-�$� 6�P�Z���~������� Ə����)� �2�L� V���z�������� ���%��.�H�R�� v������������� !��*�D�N�{�r��� �������޿��� &�@�J�w�nπϭϤ� ����������"�<� F�s�j�|ߩߠ߲��� �������8�B�o� f�x���������� ���4�>�k�b�t� ������������ 0:g^p�� ����	 , 6cZl���� ��/�/(/2/_/ V/h/�/�/�/�/�/�/ ?�/
?$?.?[?R?d? �?�?�?�?�?�?�?�? O O*OWONO`O�O�O �O�O�O�O�O�O__ &_S_J_\_�_�_�_�_ �_�_�_�_�_o"oOo FoXo�o|o�o�o�o�o �o�o�oKBT �x������ ���G�>�P�}�t� ������������� �C�:�L�y�p����� �����ܟ���?� 6�H�u�l�~������� �د���;�2�D� q�h�z�������ݿԿ � �
�7�.�@�m�d� vϣϚϬ��������� �3�*�<�i�`�rߟ� �ߨ����������/� &�8�e�\�n���� ����������+�"�4� a�X�j����������� ������'0]T f������� �#,YPb� �������/ /(/U/L/^/�/�/�/ �/�/�/�/�/??$? Q?H?Z?�?~?�?�?�? �?�?�?OO OMODO VO�OzO�O�O�O�O�O �O_
__I_@_R__ v_�_�_�_�_�_�_o ooEo<oNo{oro�o �o�o�o�o�o A8Jwn��� ������=�4��F�s�j�|�����̍�  H55�1���2�R78�2�50�J61�4�ATUP�5�45�6�VCA�M�CUIF�2�8H�NRE�52�;�R63�SCH��DOCV��CS]U�869�0��EIOCl�4��R{69;�ESET$�v:�J7:�R68��MASK�PRXuYT�7�OCO�3$������37�J�6
�53��He�L{CH�OPLG$��0O�MHCR �SMATk�MCS�#�0��55�MD�SW�B�OPB�M�PRC���s�0�PCMS�5J�������s�51/�51{�0n/�PRS�697��FRDG�FREQn�MCN�93��SNBAx�f�SH�LB�M
ǀ���2��HTC#�TMI�L􈳖TPA˖T7PTX<�EL۶��ⳗ8�����J95�_�TUTC�UEV��UEC�UFR�G�VCC��OǦV�IPG�CSCk�C�SGk���I�WE�B#�HTT#�R6lv���CG6�IG�oIPGS\�RCGƻDGB�H75/�Ru7�Ry�R66O��2O�R6�R55���4��5��D06:�F�CLI3�.��CMS˖0�#�ST-Y��TO7�7��t��_�ORSǦ��Mn��NOM˖OL��$���OPIs�SE�ND�L��Sy�EcTSsּ�S�CPk�wFVR˖IPNG�Gene�È6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p������	  H�551��2�
R�782�50�	J�614�	ATUP�5456�	V�CAM�	CUIFv28lNRE�
�52[R63�S{CH�	DOCV�wCSU�
869�0+EIOC�4�R69[ESE�T<ZJ7ZR6�8�
MASK�	P�RXY|7�
OC�OL,3<X 3��*J653�H��,LCH�*OPL�G<0�*MHCR��*SJ;MAT�MkCS;0[+55+�MDSW�;�+OP��+MPR�*��,0.PCM{5KX �+X0�+51K51�[L0KPRSK+6�9�*FRDkFR�EQ�
MCN�
9=3SNBA��+/SHLB�JM[���<2HTC;T�MIL��TPA�*TPTX\ZEL��JX0�8
�
J�95�TUT�*U�EVK*UEC�*U�FRkVCC+lO�k:VIPkZCSCN�ZCSG��I�	wWEB;HTT;�R6��\CG�kI�G�kIPGS�jR�CkZDG�+H75�KR7:+RYLR6�6�,2�*R6�R�55k|4�[5�{D�06+F�|CLI�<JCMS*�p;�STY[kTO�k78���ORSk:x �M�LNOM*OqL�;�0�OPI�j�SEND�
L:kS�Y�ETS�j {[C�P�FVR*IP=NkZGene�� R�d�v���������П �����*�<�N�`� r���������̯ޯ� ��&�8�J�\�n��� ������ȿڿ���� "�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZl~� ������  2DVhz��� ����
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �$�6�H�Z�l�~��� ����Ɵ؟���� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п �����*�<�N�`� rτϖϨϺ������� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� ������,>P�bt������� STD�LANG��	 '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�Z�RBT�OPTN�_�_�_�_�_DPN�oo*o<oNo `oro�o�o�o�o�o�o��oted ��>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� ���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _*_<_N_`_r_�_�_ �_�_�_�_�_oo&o 8oJo\ono�o�o�o�o �o�o�o�o"4F Xj|����������0�B�  �K�i�{�������Í�99ʅ�$FE�AT_ADD ?_	�������?  	ǈ� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O��O�DEMO �Y��    ǈ1]'_9_f_]_o_�_ �_�_�_�_�_�_�_,o #o5oboYoko�o�o�o �o�o�o�o�o(1 ^Ug����� ���$��-�Z�Q� c�������Ə��Ϗ� � ��)�V�M�_��� ������˟��� �%�R�I�[������ ����ǯ����!� N�E�W���{������� ÿݿ����J�A� Sπ�wω϶ϭϿ��� �����F�=�O�|� s߅߲ߩ߻������ ��B�9�K�x�o�� ������������ >�5�G�t�k�}����� ��������:1 Cpgy���� � �	6-?l cu������ �/2/)/;/h/_/q/ �/�/�/�/�/�/�/? .?%?7?d?[?m?�?�? �?�?�?�?�?�?*O!O 3O`OWOiO�O�O�O�O �O�O�O�O&__/_\_ S_e_�_�_�_�_�_�_ �_�_"oo+oXoOoao �o�o�o�o�o�o�o�o 'TK]�� �������� #�P�G�Y���}����� ����׏����L� C�U���y�������ܟ ӟ��	��H�?�Q� ~�u�������دϯ� ���D�;�M�z�q� ������Կ˿ݿ
�� �@�7�I�v�m�ϙ� ������������<� 3�E�r�i�{ߕߟ��� ��������8�/�A� n�e�w�������� �����4�+�=�j�a� s��������������� 0'9f]o� �������, #5bYk��� �����(//1/ ^/U/g/�/�/�/�/�/ �/�/�/$??-?Z?Q? c?}?�?�?�?�?�?�? �? OO)OVOMO_OyO �O�O�O�O�O�O�O_ _%_R_I_[_u__�_ �_�_�_�_�_oo!o NoEoWoqo{o�o�o�o �o�o�oJA Smw����� ����F�=�O�i� s�������֏͏ߏ� ��B�9�K�e�o��� ����ҟɟ۟���� >�5�G�a�k������� ίůׯ����:�1� C�]�g�������ʿ�� ӿ ���	�6�-�?�Y� cϐχϙ��Ͻ����� ���2�)�;�U�_ߌ� �ߕ��߹�������� .�%�7�Q�[���� �����������*�!� 3�M�W���{������� ��������&/I S�w����� ��"+EO| s������� //'/A/K/x/o/�/ �/�/�/�/�/�/?? #?=?G?t?k?}?�?�? �?�?�?�?OOO9O COpOgOyO�O�O�O�O �O�O_	__5_?_l_ c_u_�_�_�_�_�_�_ ooo1o;oho_oqo �o�o�o�o�o�o
 -7d[m�� �������)� 3�`�W�i�������̏ ÏՏ����%�/�\� S�e�������ȟ��џ �����!�+�X�O�a� ������į��ͯ��� ��'�T�K�]����� ������ɿ������ #�P�G�Yφ�}Ϗϼ����������  �+�=�O�a�s� �ߗߩ߻�������� �'�9�K�]�o��� ������������#� 5�G�Y�k�}������� ��������1C Ugy����� ��	-?Qc u������� //)/;/M/_/q/�/ �/�/�/�/�/�/?? %?7?I?[?m??�?�? �?�?�?�?�?O!O3O EOWOiO{O�O�O�O�O �O�O�O__/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O_Y  XQ/_ A_S_e_w_�_�_�_�_ �_�_�_oo+o=oOo aoso�o�o�o�o�o�o �o'9K]o �������� �#�5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ����)�;�M�_� q���������˿ݿ� ��%�7�I�[�m�� �ϣϵ���������� !�3�E�W�i�{ߍߟ� ������������/� A�S�e�w����� ��������+�=�O� a�s������������� ��'9K]o �������� #5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� ����������/ ASew���� ���+=O as������ �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? �?�?�?�?�?�?OO 1OCOUOgOyO�O�O�O@�O�O�O�O	_QPX3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u��������� Ͽ����)�;�M� _�qσϕϧϹ����� ����%�7�I�[�m� ߑߣߵ��������� �!�3�E�W�i�{�� ������������� /�A�S�e�w������� ��������+= Oas����� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�? �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o !3EWi{� �������� /�A�S�e�w������� ��я�����+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ� ���#�5�G�Y�k�}� ������ſ׿���� �1�C�U�g�yϋϝπ����������	����$FEAT_DEMOIN   ԫ�K�� �3�I�NDEX@�Oш�3�ILECOMP Z������N�.�w�SETUP2 [������  N� ��t�_AP2B�CK 1\�� � �)�����%��� ����H�� ��t���'����]� ����(���L���p� �����5�����k�  ��$��1Z��~ ��C�g�� 2�Vh��� ?��u
/�./@/ �d/��/�/)/�/M/ �/�/�/?�/<?�/I? r??�?%?�?�?[?�? ?O&O�?JO�?nO�O O�O3O�OWO�O�O�O "_�OF_X_�O|__�_ �_A_�_e_�_o�_0o �_To�_ao�oo�o=o �o�oso�o,>�o b�o��'�K��o������P��� 2��*.VR�g��p*j����s0�����uQ�PC�>�pFR6:֏���;�ʋT_�_�q�� �\���B�,����vG*.FT���q	�������C�қSTM c�l�w��d�����piPend�ant Pane	l��қH�������p��3�L�ӚGIFV������l�)�;�пӚJPGڿϋ�𿭿���T�ˊJS^χ��p��u�2�%
JavaScript��޿CS��ߊ��ϵ�� %Casca�ding Sty�le Sheet�s7ߩp
ARGN?AME.DTf��|��\z�8ߚ��Ի��g���DISP* �ߔߎ���>���0�?����	PANEL15��%�����ﵯǯu�2����������o�z�3;������L�^���z�4��%�������wr�TPEINS.XML~��:\�PbCu�stom Too�lbar���PA?SSWORDC�~?FRS:\�� %Passw�ord ConfCigW��4�/�� �[U�/qֱ䘯� ��/�b_/v���/%J(�/g/y/?'2T/=?H(+?�/�/�? ��?�/U5�?o?�?O'3\?EOH(3O�?O �O���O�?]E�OwO�O_'4dOM_H(;_�O _�_�_�OeU�__ �_&o�Jo�no�� �o3o�oWo�o�o�o" �oFX�o|�� A�e���0�� T��M������=�ҏ �s����,�>�͏b� 񏆟�'���K���o� ٟ���:�ɟ^�p��� ��#���ʯY��}�� ����H�ׯl���e��� 1�ƿU������ ϯ� D�V��z�	Ϟ�-�?� ��c��χ���.߽�R� ��v߈�߬�;����� q���*����`��� ���}��I���m�� ���8���\�n���� !���E�W���{��� 	F��j����/ �S����B ��x�+���a�,�$FIL�E_DGBCK �1\������ < ��)
SUMMA�RY.DG/�]M�D::/z/�D�iag Summ�ary{/([CONSLOGp/S/e!�/��/�!Conso?le log�/�\?TPACCN�/Y?�%A?~?�%TP �Accounti�n ?�Y@6:IP�KDMP.ZIP��?�
�?O�%�0E�xception�O�*�_\O��bQJO�_1FR DT Files�O��<f MEMCHECCKt?�/i/_1�Memory D�ata_�
l?�)	FTP�/f_��Oj_W1mme�`TBD�_�L �>I)ETHERNET�_��A�_�o�!Ether�net 0fig�ura&O�}QDCSVRF�_m__�o�Q%]` ve�rify all��o�M.cXeDIFF�ovo�o P�%�hdiff��g�A]`CHG01�o��a5��b- `y2�� &�1��gr3����� <�я`��VTRNDIAG.LS֏����.�z!Q� Ope>c� Log �!no�stic���)VDEV�DA}O�����a�VisQ�DevisceX�e�IMG��?����4�7�ʔI�mag֟c�UP�{�ESz��FR�S:\z��O@Up�dates Li�st���"�FL?EXEVENo��%�>��a� UI�F Ev�QU�?� � ,�sz)
P�SRBWLD.C	Mj��������0�PS_ROBOW�EL�_�*�HADOW4��+�D�S�Shadow �Chang�O���a��RCME�RR<�!�3���S���CFG Err{orАtailkϟ =��B��SGLIB�ϧϹ�N�:!Q� St?`_������):�Z�DU_��7���WZMDT�adn����NOTIbo�߽�R��UNotifiqc?b��t��AGXbGIGE��/�A���]�GigEZ�d��N�A��-��Q� �^������:����� p���);��_�� ��$�H�l� �7�[m��  ��V�z/!/ �E/�i/�v/�/./ �/R/�/�/�/?�/A? S?�/w??�?�?<?�? `?�?�?O+O�?OO�? sO�OO�O8O�O�OnO _�O'_9_�O]_�O�_ _�_�_F_�_j_�_o �_5o�_Yoko�_�oo �o�oTo�oxo�o C�og�o��,� P�����?�Q� �u����(���Ϗ^� 󏂏�)���M�܏q� �����6�˟ݟl�� ��%���2�[���� ����D�ٯh������ 3�¯W�i�������� @����v�Ϛ�/�A� пe����ϛ�*Ͽ�N� ���τ�ߨ�=���J� s�ߗ�&߻���\��� ���'��K���o�� ��4���X������ #���G�Y���}���� ��B���f�����1 ��U��b��>���t	�$F�ILE_FRSP�RT  ���� ����$MDONLY �1\8�  
 ��{���� ����///�S/ �w/�//�/</�/�/ r/?�/+?�/8?a?�/ �??�?�?J?�?n?O O�?9O�?]OoO�?�O "O�OFO�O�O|O_�O 5_G_�Ok_�O�_�_0_ �_T_�_�_�_o�_Co��_Poyo"VISB�CKV@e*.�VD�o�o8`FR�:\�`ION\DOATA\�oZb8`�Vision VD file�o o>Pfot^o�' ��]���(�� L��p�����5�ʏ ܏�� ���$���5�Z� �~������C�؟g� ������2���V�h�#� �����?����u�
� ��.�@�ϯd�󯈿��)���LUI_C�ONFIG ]�8�aɻ $ ��[{8 �2��D�V�h�zψ��|x ������������
ܠ� -�?�Q�c�u�߆߫� �������ߊ��)�;� M�_�q������� ������%�7�I�[� m�������������� ��!3EWi  ������~ /ASe��� ���h�//+/ =/O/�s/�/�/�/�/ �/d/�/??'?9?K? �/o?�?�?�?�?�?`? �?�?O#O5OGO�?kO }O�O�O�O�O\O�O�O __1_C_�Og_y_�_ �_�_�_X_�_�_	oo -o�_>ocouo�o�o�o Bo�o�o�o)�o M_q���>� ����%��I�[� m������:�Ǐُ� ���!���E�W�i�{� ����6�ß՟���� ���A�S�e�w��� � ����ѯ������+� =�O�a�s�������� Ϳ߿�Ϛ�'�9�K� ]�oρ�ϥϷ����� ���ϖ�#�5�G�Y�k� }�ߡ߳��������� ���1�C�U�g�y�	����x����$F�LUI_DATA ^�������R�ESULT 2_����� �T��/wizar�d/guided�/steps/Expert��"�4� F�X�j�|���������������Cont�inue wit�h G��ance ��1CUgy�`����� ���-����0 �������$���ps�o��� �����/#/5/ ���\/n/�/�/�/�/ �/�/�/�/?"?4?F>�$(:Jrip�X�?�?�?�?O O*O<ONO`OrO�OC/ �O�O�O�O�O__&_ 8_J_\_n_�_�_Q?c?ȭ_�?EJ�Ti�meUS/DST �_"o4oFoXojo|o�o�o�o�o�o��Enabl
.@ Rdv�����
��� �_��_�_f24or����� ����̏ޏ����&� �o�o\�n��������� ȟڟ����"�4�����)�;�M�zon 
`7�ʯܯ� ��$��6�H�Z�l�~���E�ST Ea�rn? Stand���� ��ӿ���	��-�?�`Q�c�uχ�� ���t�f�x�:���acces�?�+�=� O�a�s߅ߗߩ߻��������nect �to Network���%�7�I�[� m���������ȅ�A��Ϻ��ϊ�!���`Introd?uction��t� �������������� (�OL^p�� ����� $5�_�P*����V?Editor5� ���
//./@/R/�d/v/5 Touc�h Panel �� (recommen�P)�/�/�/ �/�/?#?5?G?Y?k?}?�̬P�^�?�B �?OO/OAOSOeOwO �O�O�O�O�O<�O_ _+_=_O_a_s_�_�_�_�_�_�Y�0�?�:�?o�?EoWoio{o �o�o�o�o�o�o�o �OASew�� �������+� �_�_op�2o������ ͏ߏ���'�9�K� ]�o�.������ɟ۟ ����#�5�G�Y�k� }�<���`�¯����� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ���ώ��ϲ��֯;� M�_�q߃ߕߧ߹��� ������%��I�[� m����������� ���!���B��f�(� *������������� /ASew6� �����+ =Oas2��V�� ���//'/9/K/ ]/o/�/�/�/�/�/� �/�/?#?5?G?Y?k? }?�?�?�?�?��� �?O�COUOgOyO�O �O�O�O�O�O�O	__ �/?_Q_c_u_�_�_�_ �_�_�_�_oo�? O �?Dono0O�o�o�o�o �o�o%7I[ m,_������ ��!�3�E�W�i�(o :oLo^o���o���� �/�A�S�e�w����� ����~�����+� =�O�a�s��������� ͯ�������ԏ9�K� ]�o���������ɿۿ ����П5�G�Y�k� }Ϗϡϳ��������� ��ޯ��d�&��� �߯���������	�� -�?�Q�c�"�t��� ����������)�;� M�_�q�0ߒ�T߶�x� ����%7I[ m������� �!3EWi{ ���������/ ��//A/S/e/w/�/�/ �/�/�/�/�/??� =?O?a?s?�?�?�?�? �?�?�?OO�6O� ZO/O�O�O�O�O�O �O�O_#_5_G_Y_k_ *?�_�_�_�_�_�_�_ oo1oCoUogo&O�o JO�o�o�_�o�o	 -?Qcu��� �|_����)�;� M�_�q���������xo �o�o���o7�I�[� m��������ǟٟ� ����3�E�W�i�{� ������ïկ���� ʏ��8�b�$����� ����ѿ�����+� =�O�a� ��ϗϩϻ� ��������'�9�K� ]��.�@�R���v��� �����#�5�G�Y�k� }����r������� ��1�C�U�g�y��� �������ߒߤ��� -?Qcu��� ������); M_q����� ��//������X/ /�/�/�/�/�/�/ �/?!?3?E?W?h? �?�?�?�?�?�?�?O O/OAOSOeO$/�OH/ �Ol/�O�O�O__+_ =_O_a_s_�_�_�_�_ �O�_�_oo'o9oKo ]ooo�o�o�o�ovO�o �O�o�O#5GYk }������� ��_1�C�U�g�y��� ������ӏ���	��o *��oN�������� ��ϟ����)�;� M�_����������˯ ݯ���%�7�I�[� �|�>�����v�ٿ� ���!�3�E�W�i�{� �ϟϱ�p�������� �/�A�S�e�w߉ߛ� ��l��������ƿ+� =�O�a�s����� ���������'�9�K� ]�o������������� ���������,V� }������� 1CU�y� ������	// -/?/Q/"4F�/ j�/�/�/??)?;? M?_?q?�?�?�?f�? �?�?OO%O7OIO[O mOO�O�O�Ot/�/�/ �O�/!_3_E_W_i_{_ �_�_�_�_�_�_�_�? o/oAoSoeowo�o�o �o�o�o�o�o�O�O �OL_s���� �����'�9�K� 
o\���������ɏۏ ����#�5�G�Y� z�<��`şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� j�̿��𿲟�)�;� M�_�qσϕϧϹ��� �������%�7�I�[� m�ߑߣߵ������� �߼���B���{� ������������� �/�A�S��w����� ����������+ =O�p2��j� ���'9K ]o���d��� ��/#/5/G/Y/k/ }/�/�/`���/�/ �?1?C?U?g?y?�? �?�?�?�?�?�?�O -O?OQOcOuO�O�O�O �O�O�O�O�/�/�/ _ J_?q_�_�_�_�_�_ �_�_oo%o7oIoO moo�o�o�o�o�o�o �o!3E__(_ :_�^_����� �/�A�S�e�w����� Zo��я�����+� =�O�a�s�������h z��'�9�K� ]�o���������ɯۯ ���#�5�G�Y�k� }�������ſ׿��� ��̟ޟ@��g�yϋ� �ϯ���������	�� -�?���P�u߇ߙ߫� ����������)�;� M��n�0ϒ�TϹ��� ������%�7�I�[� m�������������� ��!3EWi{ ��^������� /ASew�� �������/+/ =/O/a/s/�/�/�/�/ �/�/�/�?�6?� �/o?�?�?�?�?�?�? �?�?O#O5OGO/kO }O�O�O�O�O�O�O�O __1_C_?d_&?�_ �_^O�_�_�_�_	oo -o?oQocouo�o�oXO �o�o�o�o); M_q��T_�_x_ ���_�%�7�I�[� m��������Ǐُ� �o�!�3�E�W�i�{� ������ß՟矦� ��>� �e�w����� ����ѯ�����+� =���a�s��������� Ϳ߿���'�9��� 
��.���R������� �����#�5�G�Y�k� }ߏ�N����������� ��1�C�U�g�y�� ��\�nπ����	�� -�?�Q�c�u������� ��������); M_q����� ��������4��[ m������ �/!/3/��D/i/{/ �/�/�/�/�/�/�/? ?/?A? b?$�?H �?�?�?�?�?OO+O =OOOaOsO�O�O�?�O �O�O�O__'_9_K_ ]_o_�_�_R?�_v?�_ �?�_o#o5oGoYoko }o�o�o�o�o�o�o�O 1CUgy� ������_��_ *��_�c�u������� ��Ϗ����)�;� �o_�q���������˟ ݟ���%�7��X� �|���R���ǯٯ� ���!�3�E�W�i�{� ��L���ÿտ���� �/�A�S�e�wω�H� ��l����Ϣ���+� =�O�a�s߅ߗߩ߻� ���ߞ���'�9�K� ]�o��������� ���Ͼ��2���Y�k� }��������������� 1��Ugy� ������	 -�����"��F�� ����//)/;/ M/_/q/�/B�/�/�/ �/�/??%?7?I?[? m??�?Pbt�?� �?O!O3OEOWOiO{O �O�O�O�O�O�/�O_ _/_A_S_e_w_�_�_ �_�_�_�_�?�?�?(o �?Ooaoso�o�o�o�o �o�o�o'�O8 ]o������ ���#�5��_V�o z�<o����ŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u���F��� j�̯�����)�;� M�_�q���������˿ ݿ����%�7�I�[� m�ϑϣϵ����Ϙ� �ϼ�����W�i�{� �ߟ߱���������� �/��S�e�w��� �����������+� ��L��p���F���� ������'9K ]o�@���� ��#5GYk }<���`������ //1/C/U/g/y/�/ �/�/�/�/��/	?? -???Q?c?u?�?�?�? �?�?����?&O� MO_OqO�O�O�O�O�O �O�O__%_�/I_[_ m__�_�_�_�_�_�_ �_o!o�?�?OOxo :O�o�o�o�o�o�o /ASew6_� �������+� =�O�a�s���DoVoho ʏ�o���'�9�K� ]�o���������ɟ� ����#�5�G�Y�k� }�������ůׯ���� ���ޏC�U�g�y��� ������ӿ���	�� ڟ,�Q�c�uχϙϫ� ����������)�� J��n�0��ߧ߹��� ������%�7�I�[� m��ߣ�������� ���!�3�E�W�i�{� :ߜ�^��������� /ASew�� ������+ =Oas���� ������/���K/ ]/o/�/�/�/�/�/�/ �/�/?#?�G?Y?k? }?�?�?�?�?�?�?�? OO�@O/dOvO:? �O�O�O�O�O�O	__ -_?_Q_c_u_4?�_�_ �_�_�_�_oo)o;o Mo_oqo0OzOTO�o�o �O�o%7I[ m�����_� ��!�3�E�W�i�{� ������Ï�o�o�o�� ��oA�S�e�w����� ����џ������ =�O�a�s��������� ͯ߯���ԏ��� 
�l�.�������ɿۿ ����#�5�G�Y�k� *��ϡϳ��������� ��1�C�U�g�y�8� J�\��߀�����	�� -�?�Q�c�u���� ��|�������)�;� M�_�q����������� �ߜ߮���7I[ m������ ��� EWi{ �������/ /��>/ b/$�/�/ �/�/�/�/�/??+? =?O?a?s?�/�?�?�? �?�?�?OO'O9OKO ]OoO./�OR/�Ov/�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�?�_�_ oo1oCoUogoyo�o �o�o�o�O�o�O�O �o?Qcu��� �������_;� M�_�q���������ˏ ݏ����o4��oX� j�.�������ǟٟ� ���!�3�E�W�i�(� ������ïկ���� �/�A�S�e�$�n�H� ����~������+� =�O�a�sυϗϩϻ� z�������'�9�K� ]�o߁ߓߥ߷�v��� �����п5�G�Y�k� }������������ ���1�C�U�g�y��� ������������	�� ������`"��� ����); M_������ ��//%/7/I/[/ m/,>P�/t�/�/ �/?!?3?E?W?i?{? �?�?�?p�?�?�?O O/OAOSOeOwO�O�O �O�O~/�/�/_�/+_ =_O_a_s_�_�_�_�_ �_�_�_o�?o9oKo ]ooo�o�o�o�o�o�o �o�o�O2�OV_ }������� ��1�C�U�g�x�� ������ӏ���	�� -�?�Q�c�"��F�� jϟ����)�;� M�_�q���������x� ݯ���%�7�I�[� m��������t�ֿ�� ������3�E�W�i�{� �ϟϱ���������� ʯ/�A�S�e�w߉ߛ� �߿��������ƿ(� �L�^�"߅���� ��������'�9�K� ]�߁����������� ����#5GY� b�<��r���� 1CUgy� ��n����	// -/?/Q/c/u/�/�/�/ j���/?�)?;? M?_?q?�?�?�?�?�? �?�?O�%O7OIO[O mOO�O�O�O�O�O�O �O�/�/�/�/T_?{_ �_�_�_�_�_�_�_o o/oAoSoOwo�o�o �o�o�o�o�o+ =Oa _2_D_�h_ �����'�9�K� ]�o�������doɏۏ ����#�5�G�Y�k� }�������r���� ��1�C�U�g�y��� ������ӯ������ -�?�Q�c�u������� ��Ͽ���ğ&�� J��qσϕϧϹ��� ������%�7�I�[� l�ߑߣߵ������� ���!�3�E�W��x� :Ϝ�^���������� �/�A�S�e�w����� ��l�������+ =Oas���h� ������'9K ]o������ ����#/5/G/Y/k/ }/�/�/�/�/�/�/�/ �?�@?R?/y?�? �?�?�?�?�?�?	OO -O?OQO/uO�O�O�O �O�O�O�O__)_;_ M_?V?0?z_�_f?�_ �_�_oo%o7oIo[o moo�o�obO�o�o�o �o!3EWi{ ��^_�_�_���_ �/�A�S�e�w����� ����я����o�+� =�O�a�s��������� ͟ߟ����H� 
�o���������ɯۯ ����#�5�G��k� }�������ſ׿��� ��1�C�U��&�8� ��\���������	�� -�?�Q�c�u߇ߙ�X� ����������)�;� M�_�q����f�x� ������%�7�I�[� m�������������� ����!3EWi{ ��������� ��> �ew�� �����//+/ =/O/`s/�/�/�/�/ �/�/�/??'?9?K? 
l?.�?R�?�?�? �?�?O#O5OGOYOkO }O�O�O`/�O�O�O�O __1_C_U_g_y_�_ �_\?�_�?�_�?�_o -o?oQocouo�o�o�o �o�o�o�o�O); M_q����� ���_��_4�F�
 m��������Ǐُ� ���!�3�E�i�{� ������ß՟���� �/�A� �J�$�n��� Z���ѯ�����+� =�O�a�s�����V��� Ϳ߿���'�9�K� ]�oρϓ�R���v��� �Ϭ��#�5�G�Y�k� }ߏߡ߳������ߨ� ��1�C�U�g�y�� ���������϶��� ��<���c�u������� ��������); ��_q����� ��%7I� �,��P����� �/!/3/E/W/i/{/ �/L�/�/�/�/�/? ?/?A?S?e?w?�?�? Zl~�?�OO+O =OOOaOsO�O�O�O�O �O�O�/�O_'_9_K_ ]_o_�_�_�_�_�_�_ �_�?o�?2o�?Yoko }o�o�o�o�o�o�o�o 1CTogy� ������	�� -�?��_`�"o��Fo�� ��Ϗ����)�;� M�_�q�����T��˟ ݟ���%�7�I�[� m����P���t�֯�� ���!�3�E�W�i�{� ������ÿտ翦�� �/�A�S�e�wωϛ� �Ͽ����Ϣ��Ư(� :���a�s߅ߗߩ߻� ��������'�9��� ]�o��������� �����#�5���>�� b���N߳��������� 1CUgy� J�����	 -?Qcu�F��� j�����//)/;/ M/_/q/�/�/�/�/�/ �/�??%?7?I?[? m??�?�?�?�?�?� ���0O�WOiO{O �O�O�O�O�O�O�O_ _/_�/S_e_w_�_�_ �_�_�_�_�_oo+o =o�?O O�oDO�o�o �o�o�o'9K ]o�@_���� ���#�5�G�Y�k��}���No`oroԏ���$FMR2_GR�P 1`���� �C4�  B��p	 �p�0��F@ F�E��Q�F����C��L�FZ!�D�`�D�� �BT��@���^�?�  ������6������5�Zf5�ES<Α^�A�  ����BH��\��@�3�3@�� ����@�Q��@�g�]��Q����<�z�<��ڔ=7�<��
;;�*�<���^�8ۧ��9k'V8���8���7ג	8(��~������=�(�a�L����w�_�CFG a�T�0���ӿ�����NO� �
F0�+� 0���RM_C�HKTYP  ��p	�����RO=MF�_MINL��sW��x��7�X��SSB��b�� ��ϙu�����ϝ�TP_D�EF_OW  �t	���IRCO�MK����$GENOVRD_DOmƹ�q*�THRm� �dG�d0�_ENB�� 0�RAVC���c���� �@>�����v���^�����.� ��OU*��i�3�.��.�<u�����,��z����sC�  AD����l��$�@��B�/��1�m���.��SMT��j���������$HOST�C��1k���й�� MC�t�����v  �27.0 1��  e��BTfx �
0�������	anonymous4FXj |�r������� ��)
//./@/R/ �v/�/�/�/�i/ �/??*?<?N?�� ��?�/�?��?�?O O�/�?JO\OnO�O�? �O�/�O�O�O�O_S? �Ow?�?j_�O�?�_�_ �_�_�_+Ooo0oBo Tow_�O�O�o�o�o�o �o'_9_K_]__o5�_ t�����_�� ��(�K}o�op��� �������o13� $�gH�Z�l�~���� ��Ɵ؟����Q�� D�V�h�z���Ϗ�� �����;��.�@�R� d������������� %���*�<�N�`ϣ� ��ǯ��ۿ������ �&�i�J�\�n߀ߒ� ��7����������"��o���ENT 1l~���  P!��.s�  u�a�� ��������
���� ��?�d�'���K���o� ����������*��N r5�Yk�� ���8�1n ]�U�y��� �/4/�X//|/?/ �/c/�/�/�/�/�/?��/B?:QUIC�C0O?+?=?�?a41 �?{?�?�?a42�?�?��?>O!ROUT�ER?OO-O�O!�PCJOG�OjO�!192.16?8.0.10h?]3?CAMPRT�O�O�!�E1�@_�FR�TXO
__}_C�NA�ME !P�!�ROBO�O�_S_�CFG 1kP�� �Au�to-start{ed��FTP��a�Ϧ�Ao��eowo �o�o�oF��o�o�o *o�oOas�� �r��_oo�'Io �<�N�`�r�5���� ��̏ޏ����&�8� J�\�n�g�yϋϝ�� ������"�4�F�	� j�|�������՟W�� ����0�B������� �������ҿ���� �ݯ>�P�b�tφϩ� +ϼ���������Y� k�}�/ߑς�ſ�߸� �����߱��$�6�H� k�l��ߐ������� ��-�?�Q�2�e�V��� z�������s������� 
?���;dv� ������%�9 [�<N`r�G� �����&/8/ J/\/n/�/���� ��//?"?4?F?X? /|?�?�?�?�?�/i?��?OO0OBOTO�Z_?ERR m�Z\O�lFPDUSIZ � �0^0��D�>�EWRD ?��U�!�  ?guest�6�O��O __$_6_�TSC�D_GROUP [3n�\ �Q�9wIFT|^$PA|^wOMP|^ |^�_SH|^ED�_ �$C|^COMn@T�TP_AUTH �1o{K <!iPendanBW�Mn�[�2�q!K?AREL:*MoVohmKC}o�o�ou`�VISION �SETfP�o�o�v! ,rcP>hb�������~dC�TRL p{M�6��1
F�FF�F9E3��$F�RS:DEFAU�LT[�FAN�UC Web Server[�I��" d�O�D�я������+�jDWR_CONFIG qkU��Bc[�lAI�DL_CPU_P5Cz��1B�� ��w BH��MIN���sQ��GNR_IO�uA�B�0�H��NPT_SIM_DOӖ�ݛSTAL_S�CRNӖ �ޚT�PMODNTOL8�ݛ��RTY�������` `ENB��sS��OLNK 1r{KxP����ɯۯ�������MAST�EҐy�5���SL�AVE s{KH� D��SRAMC�ACHE/�A�"aO�_CFGq�����U�O�`����CMT_�OPz�ՒJǳYC�Lp���t�_ASG� 1t`��A
  �6�H�Z�l�~ϐϢ� ����������� ���	�NUM�CI
慲IPn���RTR�Y_CNҿ���_�UP_��A����E ؅�����u)�  �06��م�RCA_ACC 2vk[�  R�� ��i � 5� 7Þ�0�i��,�. s p#��  �2�D���BUF001� 2wk[= {�u��u0��������#��2��C��Vu0�% Pou0�Bx2��u0��q�������u0�sP����Ц��������"�  "�ۋJ��U.�cu�0�r`�|u0Z�p��.�U�.��.��.��.���.�Ԗ�So2��  2�S�~���u0!�SpS��u0X]�S��~��~��u0��p�S���T�q  �qT ���/��@��d� _ �Tz�����������R���������R��=��r�䃲�䒖�]�������s�2���d���������� ����������t� ���tp =���t� x�� ����������%�&�,�``�4��<�AE� AM�AU�A]�Ae� Am�Au�A}���<���e �� ���������������������W������������U (�����kX	�" � � ���	l�,>Pbt003 ��� ���1�� �"����"����"�� �"��"����"��" ��"�#�"%�3 :25�C:2E�:2M�[ :2]�k:2m�{:2}� ��2����2��2 ���2��2����2 �������2����2 ��#�#�"## �"�$5#� �$E#� O4 U#� ^"� f"� o4u#`� ~"���я�2xk[G 46�A��Q�P�<�P�D�AՒ��H�IS}�zk[ ��� 2021-�04-21�V � ;qb'_9_ K_]_o_�_�_�_�_�_� L[T�Q18?-02-27Y�_�
oo.o��T�8�:�PQocouo�o�o�[N���W1�A�_�o�o�\��C���BX��;W  `th&tpt�xt�&t��'s���8�9�Jo� LM���hU��o�����<��D���-r:P3ErRqt�t�tјt�2�@�t��\��RL�ڽh2� ������5�r�%r�@ -z�@=r*pEz.�@�ts��[��RK��h�Z;�z���r*pSa!'s��ҟQ���8����VJ�n�h�" a�N�`�r�r���ݍf7���ʯUQ���n�-��G� �O_Z1 sM�_�q� ��������˿ݿ��_@;�%�7�I�[�I`:�@c\χϙϫϽϫo�o ���u��Bdp=�%p�d-p=��M�=p =�Ep=��M�UpM�]p�d(ߛ߉����� ���v=������Z�t� ;��=��=��=҇� =�Q�=�Y��n����� ����ȍ��%p=�R�=� b�M�j�Q�c�u�5��� J�\�������5�Mҹ� MҼ������"4"� 4�j|�������� ��]���ާ���� �L� �&�Z�| �������/����/T/f/x/Ah �/�/�/�/�/�/��9/ &?8?J?t҅P%r� P�Pb��2"��2��3��3]p�A�?�?�� ��?OO�y7O �|; REr�3R�P�P �P%��PY��O�� �?�O�O_ʍl?ZOlO ~O�O4��_q��O�_�_ �_\?��oo�7oIo [oI[�o�o�o�_"_ �`���o�J�;��I_CFG 2�{: H
C�ycle Tim�e�aBusy>DwIdlzr�t�mi8|�q�Upvv|qRea}d�wDow8x֟ �rqsCo�unt|q	Num� qr�s�={��`��q�PROGWr-|:D�0�u����������Ϗ�y �S�DT_ISOLCw  :� ��@~J23_DSP_ENB  ��>#�INC }���e�A   ?�OP=���<#��
�j�:�o �u������a��ȟ�OBK�C,��uU���G_GROUP �1~�U�< � �j�Cy.�ПE?Dxd�m��`Q�� ����̯�����&��Dw��ڙG_IN_AUTO�Q�#��POSRE���K�ANJI_MAS�K��t�KAREL?MON :(��by���(�:�L�(@~²O��V�X���nŉ���CL_LNd�NUM0������EYLOGGIN�G��?�v�U�F�L�ANGUAGE �:
���DEFAULT l�(LGXq�V���r�4�  S8�p��`'�g'  ��`�ۏ��;��
��(U�T1:\\Ϧ�  �ߵ����������!�8�E�W��(��#�LN_DISP ��M��x������O�CTOL���aDz�@��f��GBOOK �)��z�qz�z�� 'Uy�k�}� ����������5Ӱs����	-�t�*��/�ُ`�+�_BUFF� 2�� A�Evꂒ�w �����#, YPb���������/��ZDCS �V�Y�n��� #Dx^u�/�/�/�/6$�IO 2�B+ !cp�/cp@���/? ?*?>?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO^OnO�O�O�O�%�ER_ITM��d D��O_#_5_G_Y_k_ }_�_�_�_�_�_�_�_ oo1oCoUogo	��B�SEV�����FTYP���O�o�o�o�vm��RST��4%S�CRN_FL 2��-@��g/gy������TP������b�NGN�AM,�`�
�2$UPMS��GIp��U�}B�_LOAD��G % �%D�ROP��MAXUALRM�¢� ��U�
��H�_P�RM��� !���C���7�������P 2�7� �q�	�ol�W���{� ��Ɵ���՟��� D�/�h�S�������¯ ���ɯۯ��@�+� d�v�Y����������� ��߿��<�N�1�r� ]ϖ�yϋ��Ϸ����� �&�	�J�5�n�Q�c� �ߏ��߳�������"� �F�)�;�|�g��� ������������ T�?�x�c����������������DBGDEF ��[!���_LDXDISA�-��{�#MEMO_{AP'�E ? �
 $x(�����������F�RQ_CFG ���(A x'@i�E��<[$d%�m$:������*�/� **:���� �_����+/"/4/ a/X/j/�/����/�@`�/�/�/�/�',(�/ >?�$,?i?P?�?t?�? �?�?�?�?OOOAO�(OeOwO^O�O��IS�C 1� �� � ���O��)�O��2__�V_�O�B_MSTR� ��myUSCD 1�o�N_�_J_ �_�_o�_4oo1ojo Uo�oyo�o�o�o�o�o �o0T?xc �������� �>�)�N�t�_����� ������ˏ���:� %�^�I���m������� ܟǟ ��$��H�3� l�W�i�����Ư��� կ����D�/�h�S����w�����Կj_MK�'��]Y�$M�LTARM&�:-� 3" �P�X� METPU�K ǲ���YND�SP_ADCOLxr�& }�CMNT�� ��FN���τ�FSTLI���ǁP ��^'�G�Y?�|IԆ�POSCF��=��PRPM��Y��ST��1��[ 4Q#�
��ϱ�� ���׿�������7�� +�m�O�a������ ��������E�/���SING_CHK�  ��$MODA%��K����DEV 	N
	�MC:��HSI�ZEKǰ��TA�SK %N
%$�12345678�9  2}�TRI�G 1��[ l ^9n�=�YP��5��~�E�M_INF 1���`)AT?&FV0E0�+�)E0V1&�A3&B1&D2�&S0&C1S0}=)ATZ+fH��:��bA�/�'//K/]/ �/5GYk �/� ?7/$?6?�Z? ?~?�?w?�?g/y/�? �/�/�/2O=?�/hO�? �OGOQ?�O}O�O�O
_ _�?@_�?OO)O�_ MO�_�O�_�_�Oo�_ <oNo5oro%_7_�o[_ m__�o�_&]oJ o�;���� �o��o�o�o�oX� |������e֏������0���NITO�R�G ?��  � 	EXEC�1˳s�2y�3y�4�y�5y�C {�7y�8
y�9˳t��rޔx� ޔ��ޔ��ޔ��ޔ�� ޔ��ޔ��ޔ̒ޔؒ�ޓ2�2�2��2�	�2�2!�2-�2�9�2E�2Q�3�3��3���R_GRP_SV 1� � (7�5�(�>���<����0+&��=I�?�j���
_D�ς��9�ION_D�B���Ǳ  C��~���~���Ћ����v�W�&�_N   ?��?�����̢�-ud�1����υ�PL�_NAME !�<��!De�fault Pe�rsonalit�y (from �FD)����RR2��� 1�L6��LA�<��� d:҉ϛϭϿ��� ������+�=�O�a� s߅ߗߩ߻���������2��.�@�R�d�v��������< �����0�B�T�f� x����������޲����
���P J\n���� ����"4F X'9����� ��//0/B/T/f/ x/�/�/k}�/�/�/ ??,?>?P?b?t?�?��?�?�?�?�?�> �H�6 H�b� H\���  #�O1M�dC@ PObMFO�O�G@�=��|C�O�M�O�O C �H__ _2_P_V_�t_�_�f��_�\��E	`_�_o o�Q:�oA`�@oRo�dovn A�  �i�O�o�Lޱ�o�k �O�o'9$]Ht� �R�� 1�4�����R@ �� &�<��p @D7�  �q?��s�q�?��q�A��6�Ez  �q���;��	l�r	 ��@�� 0�ް!� ���p� � �� �F��J���K ��J˷��J� �J�4�JR�<g|v�f�0O���@�S�@��;fA6A���A1UA狠X{����=��N��f������T;f���X��ڀ��*�  ��  �O5��>��p�H���?��?����#�����ԏur`�f��q{��g�������i�V�}��(  ����񤰞�ʔt柉�	�'� � ��I� �  y��e��:�È(�?È=���@������ <!��� � ��  ��qz���r�o�o����ү�  '覵��@�!�p@�a�@j��@��@��C�KC"��"��B�p�C%����@��r�  ����n�������m;a;n�`@����D�u՟ҿ �������Q�c�E��UŔ�� :�W � x�x?�ff0�O�Ϙ�*� �P����ˍ�8�����>����x��q����0�P�:�U�7�0�0���>��|���<2�!�<"7�<L���<`N<D��<��,h��ߴ��s���s ҈`?ff�f?��?&�аT@�T���?�`�?Uȩ?X� ᒩL����t,��t8� �wW�����ό�w�� ����������.��R���!�F�A��� =���)���M����HmN H[���G� F�� HZE~i��� ���� �oAK ��������)� ��/��%/7/�j/ U/�/y/�/�/��M��"�i��C�/?�/5? =8��??F??j?���ç�s��-M�BH�"��.��?,�[2�xY0X1�1@Iܔ=�@n�@���@: @l���?٧]�? ���%�n��߱���=�=�D��0OB@���@�oA�&{�C/� @�U�XO�+J8��
�H��>��=3�H��_�O �F�6�G���E�A5F�Į�E��O�@���fG��E���+E��EX���O�@>\�G��ZE�M�F�lD�
�p�O�? E_0_i_T_�_x_�_�_ �_�_�_o�_/ooSo >owobo�o�o�o�o�o �o�o=(:s ^������� � �9�$�]�H���l� ������ۏƏ���#� �G�2�W�}�h����� ş���ԟ���
�C� .�g�R���v������� �Я	���-��Q�<��u�`�r���fB(hA4g���h������3�ϩп��!�4 �{����!��0+#(�:��j�bT�f�1E���|�Ђˀ��Ϯ���P�����iP��P:�IVc߶�oߙ߄��ߨف����������9�$��"$<�N�� r�����v�H���&��e,�6�l�Z�|�����n)���������8F
  2� H�6�&H�,{�g\��&B�!�!�� B��0�0A� @ �/��$�3���l^pUgy����$0� �� ��� T�%
 ��//+/=/ O/a/s/�/�/�/�/�/��/^J� ��$�����4�$MR_�CABLE 2�>$� � V�UTP��@n�?�0�F1�?0��0z B�z C[0n�OM�`�B���n��)�� D���G??Q65  B�� T�O
�vr0���s����WD��2�貓?�7� �� C�� 9h4��r0����N~6��,�?�?�*\0�� [@�CW@j27�(Ԧn�:̉c�6E�/T3 �OR˰O�O�O�O�O_ �O�O"__*_�_�_`_ �_�_�_�_�_oAn�+��_Qocouol�?op�o�o�ol�*�o�** 3OM }�%9��zH���%% 23�45678901%7u "RFqn�[@� �n�n�
�Lw�nnot s�ent �jzsW�,�TESTFECSALGRI��gkʝd�t��q
,�tG �P�n��"���'�9�K� 9�UD1:\mai�ntenance�s.xmlS��� � ��DE�FAULT2G�RP 2�	z � pLn�  �%�1st mec�hanical �checkL}n���6��>�G�H �$r���������n���controller��7��Ic�8�J�\�n���ϑcM���n�"8��!n�ȡϯH'��� ��*�<���Cٟn�����Y����ҿ�h���ϒC�ge��. batter!yς�W�H	������ϨϺ���ϑSu�pply grecasK���È�
�!<���Hs�HߠZ�l�~ߐ�ϑ �c�abl��߾�g�
 7���0�B�T��ؑ+�����Q�����������`�$��@�hoo� ��������� ��+� O�a�s�)Z l~�����' 9 2DV� ��{����
/ /k@/R/�v/��/ �/�/�/�/1/?U/g/ <?�/`?r?�?�?�?�/ �??-?OQ?&O8OJO \OnO�?�O�?�?�OO �O�O_"_4_�OX_�O �O�_�O�_�_�_�_�_ I_om__To�_xo�o �o�o�oo�o3oEoWo >Pbt��o� �o���(�:� ��p��_����ʏ ܏� �O�$�6���Z� ��~�������Ɵ�� 9�K� �o�D�V�h�z� ��۟������5�
� �.�@�R���v�ůׯ ����п�����g� <ϋ���r����ϨϺ� ����-��Q�c�8߇� \�n߀ߒߤ������ )�;���"�4�F�X�j� �ߎ������������ ��m���T���C��� ����������3� i�>��bt��� ���/S(:�L^p��	 T ~�����// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO�fOxO  �?�  @�  ��O�O�O��O__�(_�*H_** ���@zO|_�_�_�b_�_�_�_�_�� !__�_Ko]ooo1o �o�o�ooo%o�o #5oAk}��o �oQ���E�1� C�U����a����� ӏ����	��e�w��
��$MR_HIS�T 2��v��� 
 \�$ 2�34567890�1����P�BR��9 ���������?�Q� c��,�������t��� ԯ��ί;��_�q� (���L���˿��￦� �%�ܿI� �m��6π��Z����ϐ���[�S�KCFMAP  ]�y��B�������ONREL  ���v�.�6��EXCFENB`�
,��y��FNC��r�JOG_OVLIM`�dv�\���KEY`���=��_PAN_���\���RUN�����SFSPDTYPx��k��SIGN`�>r�T1MOT��o���_CE_GRoP 1��.� ~���O��÷���a� �����C�U��y�0� ����f�������	�� -?&c��� �t�����Mq(�QZ_�EDIT]�(�Q�T�COM_CFG 1�$������� 
�_ARC_�}�`��T_MN�_MODE]�����UAP_CPL�/��NOCHEC�K ?$� �� �/�/�/�/�/ �/�/??0?B?T?f?�x?�?�?I�NO_WAIT_L\���NT��$�3�ý�1_ERR��2	�$�6ф�OEOWOiO@�L<юO�O�53 OC}�#M| �lf�³��A(C���$�8Ο,��C�#C3��r��<�� ?����_�O?�7NBPAR�AMB�$����Fg�_yW8ѫ_�[ = ���_�_�S�_o (oo4o^opoLo�o�o�kxW��o�l}_�n#UM_RSPA�CE!��b�GQt�$ODRDSP#�_��OFFSET�_CAR�_/�vDsIS��sS_A3 �ARK]�OPE?N_FILE�p_����cqPTION�_IO�����M_�PRG %3z%c$*A�S��sWO�p[����C쀸�����  ;��?֞��g��	 �h�Ȟ����4�dp�RG_DSBL  n�.�J��sRIENTTO_����C�>�-�A ��rUT_SIM_ED�+ҋBdpVhp?LCT ��=�藄O}��d\�_PEqX; ���RAT;'� d�����pUP� �m��pw����� �>�L��$P�AL�2��>`�_POS_CH�p��`��ZP2��L6��LA�W� ���oѯ�����+� =�O�a�s��������� Ϳ߿���'�9ϵ�2��h�zόϞϰ��� ������
��CW�4�F� X�j�|ߎߠ߲����� ����*
AAs'�}I5�4�Z�
BPG���� ����������&�8� J�\�n�����a�s��� ������"4FX j|������� ��0BTfx �������/0//_�xW�Y/k- ���c���/�+�/�/�'�>->-�o?�/3?�' tP(7R?H?Z?l?�?�? �?�?&0w��?L�D(4�	`<?6OHOZOA:�o<�xO�O�O�O>�`A�  �I!? �O�__�]?>_)_b_ M___�_�_�_u�����O�1������� ��$B�@ �؄��P �@D�  a?��c�Q?<�a<�D��  Ez0c�:�;��	l&b	 ��@�� 0PP_` ��
`� � �� ��b�PH0�#H��G��9G�ģG�	{Gkf���GΈK/X�o�l�PC�1��`�[�D	� D@� D7g�n�d����  �5��>�(p`�4�(: �B4�Bp{����!<���O��"��r'a�sW��Ao�Rҧpߐ}�p(  ��p�����_$��U	�'� � B��I� �  y��E�F=���f��x���� <�_`� � � ��ف��8� b__�W9N=��  'N�(�,�aOpC�`��`[pB`Cc5�G� ����@�i����m�����G�MuAuN�@@ <��*b7e����4� �X�C���������<�O� :�a�tx?�ff�/į֯�h� @��O�8x<�3�A�>�׶q"a�J�pn�Px���uaxncnd؃>�������u<2�!<"7��<L��<`N�<D��<��a,�o��c� c|^��@?fff?��?& �K�@T��2�?�`?U��?X�B�:銒 �'d�Iev�g��� Zd���ϵ�������� 6�!�Z�l�Wߐߢ�y� �߱���aσυ���D����HmN H[��ArG� F�� M���������� ���(��%�^� _� ��K�����+���g� *<N�cu@������Β���I={C�O�<s^?��}�X��?yç'c�'*sqH�`�xp�������:!@I��>}@n�@���@: @l���?٧]/ ���%�n��߱���=��=D��n/� ���@�oA��&{C/� @��U�/ �+J�8��
H��>���=3H���_�/ F�6��G��E�A5�F�ĮE����/� ��fG���E��+E���EX�?� >�\�G�ZE��M�F�lD�
`8?/�?n?�?�? �?�?�?�?O�?OIO 4OmOXO�O|O�O�O�O �O�O_�O3__W_B_ {_f_x_�_�_�_�_�_ �_oo-oSo>owobo �o�o�o�o�o�o�o =(aL�p� ������'�� K�6�H���l�����ɏ ���؏��#��G�2� k�V���z��������z�"(�!4��榱���֕3���� ��!4 �{x:�L��!�0+#f��x�Z�jb����1?E�䴛|��� �����"��F�4���%P޲Px������������׿¿��湿�� ��A�,�Q�w�bϝ"$zό��ϰ������@����@�.�d�R�ej߀tߪߘߺ�������)����.��R�@�v����  2 H��6�&H�����\�b�&B##B� 
 A� @'����� "�4�F�W���߁�@�����������$ԥ� � q�� ��%
 ��3E Wi{���������* ���b����4�$�PARAM_ME�NU ?����  �DEFPULS�E�+	WAIT�TMOUT�R�CV� SH�ELL_WRK.�$CUR_STY�L�OPT����PTB��C��R_DECSN �i�<,6/H/Z/�/~/ �/�/�/�/�/�/??� ?2?[?VSSREL_ID  ������j5USE_P�ROG %e%8W?�?k3CCR�|2���m�7_HOST7 !e!�4O��:T���?-C�?A�/CiO�;_TIME�|6�5VGDE�BUGz0ek3GI�NP_FLMSK̒O�ITR�O�GPG�A�@ �Lp� [CyH�O�HTYPEbn�V?P?�_�_�_ �_�_�_�_oo?o:o Lo^o�o�o�o�o�o�o �o�o$6_Z l~���������7��EWORD� ?	e
 	�RS�@�PNeS��s�JO!��TEP@}�CCOL�3���3WL�0� ���	���5d��ATRACECToL 1���ow v�� �������&���DT �Q���S��D� � h�t��h� n�	 �n�$Pn� n��j��*r��z���������Tn���l�l�	l�U�j��r��z����U������
l�l�l�l�k�}��������şן����� `�:�L�^�p������� ��ʯܯ&� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ�������`��
��.�@� T�QT�|0V�T�T�UT�T�T�T�UT�T�T�T�QT�! V�T�T� �Z�l�~ߐߢ�쯮� ���8�J�\�n���� \������������� "4FXj|�� �����0 BTfx���� ���//,/>/P/ b/t/�/�/�/�/�/�/ �/??(?:?L?^?p? �?�?�?�?�?�?�? O O$O6OHOZOlO~O�O �O�O�O�O�O�O_ _ 2_D_V_h_z_�_�_�_ �_���_�_
oo.o@o Rodovo�o�o�o�o�o �o�o*<N` r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P� b�t���������ο� ���_�:�L�^�p� �ϔϦϸ������� � �$�6�H�Z�l�~ߐ� �ߴ���������� � 2�D�V�h�z���� ��������
��.�@� R�d�v����������� ����*<N` r������� &8J\n� �������/�"/4/F/X)�$PG�TRACELEN�  W!  �_�V �l&�_UP ������!� �!�� l!_CFG M��%�#V!� ��$�$�/�'~ �*�  ��%�"D�EFSPD ���,U!~ �l I�N� TRL ��-�!8�%C1PE__CONFI� ��%���!�$\�)l LID�#��-�	�9LLB 1��~7 ���$B�  B4�3�& �5JO�E�/ << T!?�1KPO1OHO jO�O~O�O�O�O�O_ �O�O_L_2_T_�_�ZB�_�_�_�_3O�_�"oo'oXo�9GRP� 1��<W!@�  �[�V!�A?x�D P��DV�C2�� o�V d,D�i�i�1�0��0Wo)O�1F�n´(s
�kB+p Rq2.hR�V!�>'oY>a�����~� =N�=R��3�� 0�i�T���x����Տ�����  Dz0�9�V 
 �a��q� ��������ߟʟ�� '��$�]�H���l������)W!
V7.10beta1�$�ܠB(�A�\)A�G��a�ޡ>�������ޡA�����ffޢA�?p�AaG��Q�Q#@�(��`� ��K�0]�o����#Apأ�r �0����Ϳ߿ڢU!�� }���v�$��H�2���:KNOW_M � �%�&�4SV {��9��5N�����f�9�$ߠ6�o��"�m�3Mvc����} ��	�%���T���P��$����פ�@1ߠ���(�wPV�1MRvcĥ�T~��D��u����OAD?BANFWD�ϡ3{STva1 1ś)��4�5���� �&��� �Q�D�V�h� �������������� 
O.@�dv������2�����V �<%�w`3 !3E��4bt����5�������6//,/>/��7 [/m//�/��8�/�/X�/�/��MA���d�3�'OVLD � ;�ߊ���P�ARNUM  p��?�?��SCHS9 a5
�7�1�9��
EUPD�?�5uTO>�%_CMP_��V0�����'��lDER�_CHKzE��`��ҎFwO�KRSg����pa_MO���H_��O�%_RES_G
���;
8��oi_\_ �_�_�_�_�_�_�_o �_/o"oSoFo9?+U6\F_xo+Ua�o�o �o-S��o�o�o-S  27-SZ Rqv -S� ���-S 0�x��-RV 1���|���@`z$�BTHR_INRg��X1����dc�MASmSp� Z��MNo����MON_QUEUE ������@����$Nq@U�AN8��ۈ�END��_��EXE ��6@B�E���OPTI�O��[��PROG�RAM %Պ%��.��?�TAS�K_IU4g�OCFG �Տ�?ɟ���DATA����@(�2��k�}��� ����^�ׯ������ʯC�U�g�y�,�IN+FO���I���5� ҿ�����,�>�P� b�tφϘϪϼ����π����(�:ߕ�����I� di���@DIT ���߬���WERFLA�V����RGADJ �^��A�  ��?�@`�w����� ��W�_�?���z�N�@<@�9���%?`h���dm�C�2�%�V��	H�l7�U��2�?G�A ��t$���*��/�� **:���@�����2�5,�'�����1��1W�9�Q����/� A�o�e�w��������� ����]G=O �s����5� �'�K]� ��/����� y/#/5/c/Y/k/�/�/ �/�/�/�/Q?�/?;? 1?C?�?g?y?�?�?�? )O�?�?O	OO�O?O QOOuO�O_�O�O�O �O�Om__)_W_M___ �_�_�_�_�_�_Eo�_ o/o%o7o�o[omo�o�o�oN�	�<��* cNt����Q�M����PREF S�%�����
��?IORITY��܆}���MPDSP������C�U������OoDUCT�������OG��_T�G��钍ڂ�HIB�IT_DOA���TOENT 1Ӊ�� (!AF_�INEm� �+�!�tcp+�S�!�udB�{�!�icmj�qXY��ԉ����)�a ��ߟ����ٟ ���	�F�-�j�Q�c� ����į�������H�B�T�*����%����V����>rlD�f��/	�����һ��~��AG�,  ��o�D�V�Ph�z��պ��Z뿠�������ϻ�i�E�NHANCE )�u�s�A��d�P�7�~����������PORT_NUM�n������_CARTREP�|Ĝ�SKSTAm���SLGS���ě�G�T�Un?othingX�5��G�Y��{��TEMPG ڑ�e��e��_a_seiban���������"� �F�1�j�U���y��� ����������0 @fQ�u��� ����,P; t_������ �//:/%/^/I/[/�//�/q�VERS�IL����  disablej��m�SAVE ����	2670H�755�(�/E?!`@�G?Y?|�}? 	�8Hw��o�;�?��e�? O"O4OFOTJ�<|?�O��5_�� 1�
ě20�@r�e�Ox�O�g�pURGE�1B掘�WFP�p����W�3T�ѯ��WRUP_DEL�AY ���&UR_HOT %!v�z�?߳_DUR_NORMAL�X���_�_�WSEMI�_�_;o��qQSKIP�C�|��Cx�/�o�/�o�o �o�m}�o's�o!3 EiW���w �����/��S� A�c�������s�я�� ����ߏ�O�=�s� ����]�����˟��|�SRBTIF4T���RCVTMOU������/�DC�R�C�^i �ЗaBJ�'B��[yB��@��$�?(��)�{���mH\�e���1��p����1R�oۯ�o �<2�!<"7��<L��<`N�<D��<�� 9��O֯?�Q�@�u� ��������Ͽ�����)�;�o�RDIO�_TYPE  عM1�G�ED�T_?CFG ��Kb�BHSE��Xa2]�� �ȸ� ����.� �үD�/�h� S��ϙ�(o���o��ӟ �����;�)�_�M�� m�ߴ�9�{������ ��%��5�7�I���� ������a�������! E3i�����a �]���A /e���mG� ��/�+//O/q v/�/G/�/C/�/�/�/ �/�/'??K?m/r?�/ S?�?�?�?�?�?�?O��?!OW?}?nO;���I�NT 2�Y���_�G;� �O�K�x+��OX�f�0 _ [3O6_'OF_H_Z_�_ ~_�_�_�_�_�_o�_ 2oo*ohoVo�ozo�o �o�o�o�o
�o.@ &dR�v��� �����<�"�`��N���!�EFPOS�1 1�d�  x\O҉���O�� ��+�ŏ׏�r�]� ��1���U�ޟy�۟� ��8�ӟ\�������-� ?�y�گů����"��� F��C�|����;�Ŀ _���������B�-� f�ϊ�%Ϯ�Iϫ��� �ߣ�,���P�b��� �Iߪߕ���i��ߍ� ���L���p��� /����e�w����� 6���Z���~��{��� O���s����� 2�� ��ze�9�] ����@�d ���5G��� /�*/�N/�K/�/ /�/C/�/g/�/?�/ �/�/J?5?n?	?�?-? �?Q?�?�?�?O�?4O �?XOjOOOQO�O�O �OqO�O�O_�O_T_ �Ox__�_7_�_�_m_ _�_oo>o�_bo�_��o!o�o�oUc��2 1崏^opo�o( LRop�/�� e����6��� �/���{���O�؏s� ������2�͏V��z� ���9�K�]������ ���@�۟d���a��� 5���Y��}������ ů��`�K������C� ̿g�ɿϝ�&���J� �n�	��-�g��ϳ� �χ�߫�4���1�j� ߎ�)߲�M���q߃� ����0��T���x�� ��7����m����� ��>�������7����� ��W���{���: ��^����AS e� �$�H� li�=�a� �/���/h/S/ �/'/�/K/�/o/�/
? �/.?�/R?�/v??#? 5?o?�?�?�?�?O�? <O�?9OrOO�O1O�O�UO�O�o�d3 1� �o�O�O�OU_@_y_O �_8_�_\_�_�_�_o �_?o�_co�_o"o\o �o�o�o|o�o)�o &_�o��B� fx��%��I�� m����,���Ǐb�� �����3�Ώ���,� ��x���L�՟p����� ��/�ʟS��w���� 6�H�Z��������� =�دa���^���2��� V�߿z�Ϟ���¿�� ]�Hρ�ϥ�@���d� ���Ϛ�#߾�G���k� ��*�d��߰��߄� ��1���.�g��� &��J���n����� -��Q���u����4� ����j�������; ������4���T �x��7�[ ��>Pb� ��!/�E/�i// f/�/:/�/^/�/�/?<�OT4 1�_�/ �/?�?m?�?�/�?e? �?�?�?$O�?HO�?lO O�O+O=OOO�O�O�O _�O2_�OV_�OS_�_ '_�_K_�_o_�_�_�_ �_�_Ro=ovoo�o5o �oYo�o�o�o�o< �o`�oY�� �y��&��#�\� ������?�ȏc�u� ����"��F��j�� ��)���ğ_�蟃�� ��0�˟ݟ�)���u� ��I�үm������,� ǯP��t����3�E� W����ݿϱ�:�տ ^���[ϔ�/ϸ�S��� w� ߛϭϿ���Z�E� ~�ߢ�=���a����� �� ��D���h��� '�a�������
��� .���+�d����#��� G���k�}�����* N��r�1�� g���8?045 1�;?��1 ������/� /Q/�u//�/4/�/ X/j/|/�/??;?�/ _?�/�??�?�?T?�? x?O�?%O�?�?�?O OjO�O>O�ObO�O�O �O!_�OE_�Oi__�_ (_:_L_�_�_�_o�_ /o�_So�_Po�o$o�o Ho�olo�o�o�o�o�o O:s�2�V �����9��]� �
��V�����ۏv� ����#��� �Y��}� ���<�ş`�r����� �
�C�ޟg����&� ����\�寀�	���-� ȯگ�&���r���F� Ͽj�󿎿�)�ĿM� �q�ϕ�0�B�Tώ� ����߮�7���[��� Xߑ�,ߵ�P���t��� �ߪ߼���W�B�{�� ��:���^����������A���e�K]6 1�h�$�^�����  �$��H��E~ �=�a��� ��D/h�' �K���
/�./ �R/��/K/�/�/ �/k/�/�/?�/?N? �/r??�?1?�?U?g? y?�?O�?8O�?\O�? �OO}O�OQO�OuO�O �O"_�O�O�O_|_g_ �_;_�___�_�_�_o �_Bo�_foo�o%o7o Io�o�o�o�o,�o P�oM�!�E� i�����L�7� p����/���S���� �����6�яZ���� �S�����؟s�����  ����V��z���� 9�¯]�o������� @�ۯd�����#����� Y��}�ϡ�*�ſ׿ �#τ�oϨ�C���g� �ϋ���&���J���n��	ߒ�x���7 1� ��?�Qߋ�	���-�3� Q���u��r��F��� j������������ q�\���0���T���x� ����7��[�� ,>x���� !�E�B{� :�^����� A/,/e/ /�/$/�/H/ �/�/~/?�/+?�/O? �/�/?H?�?�?�?h? �?�?O�?OKO�?oO 
O�O.O�OROdOvO�O _�O5_�OY_�O}__ z_�_N_�_r_�_�_o �_�_�_oyodo�o8o �o\o�o�o�o�o? �oc�o�"4F� ����)��M�� J������B�ˏf�� �������I�4�m�� ��,���P���럆�� ��3�ΟW����P� ����կp�������� �S��w����6���<�߷�8 1���l� ~���6�!�Z�`�~�� ��=ϟ���s��ϗ� � ��D������=ߞ߉� ��]��߁�
���@� ��d��߈�#��G�Y� k�����*���N��� r��o���C���g��� ��������nY �-�Q�u� �4�X�|) ;u����/� B/�?/x//�/7/�/ [/�//�/�/�/>?)? b?�/�?!?�?E?�?�? {?O�?(O�?LO�?�? OEO�O�O�OeO�O�O _�O_H_�Ol__�_ +_�_O_a_s_�_o�_ 2o�_Vo�_zoowo�o Ko�ooo�o�o�o�o �ova�5�Y �}���<��`� ����1�C�}�ޏɏ ���&���J��G��� ���?�ȟc��ҿ�MASK 1����0�>��XN�O  �=�C�M�OTE  _�  ���_CFG �휭��PL_�RANG�������٦OWER ������SM_D�RYPRG %���%��I��TA�RT �	�W�U?ME_PRO&�8�����_EXEC_�ENB  ����GSPD��ΰָ;�TDB���RM��I_AIoRPUR� ���m�p��MT_�T������OBOT__ISOLC]��l��̥ȥ��NAME� �����O�B_ORD_NU�M ?	�i��H755  ���@�R�d��PC�_TIMEOUT�� x�S232浢1�`�� L�TEACH ?PENDAN�б�,С��������Mainten�ance Con%s������"�ߒ�No Use�� ���@�R�d�v������NPOf���С�����CH_�L�����	����!UD1:�1���R�VAIL�!ц�������SPACE1 2�`�
��ХЩ�刷�ΦТ�m���<o ���?�Y� Y���KlC�| ���������% <�QrY`�d�� ����Y)/ @/�U/v/]/�/�� ����//7/-?�/ Q?r?�?k?�/�/�/�/ �/�??3?)OJO	O_O �OgO�O�?�?�?�?�? OOAO7__[_|_�_ e_�O�O�O�O�O�__ =_3oToou_�oqo�o �_�_�_�_�oo)o/ Moe�]o�o�o �o�o�%G=�^� ���{������ ���!�S�9����o����g������2��� ��ݏ����%� W�Z���:�������Ưǟ3ڟ����"�ԯ F�x�{���[���ҿ����4����1�C� ��g������|��������	�5�.�@�R� d�߈ϺϽ�ߝ������)�*�6=�O�a� s߅�7������$�� �5��J�K�7^�p� ����X�������E�@��5V-kl�8� ��������y�� �f VwN��Gw �� ��ń
� �  �//1/C/U/g/ y/���-���/m�/ȁd0�/2?D? V?h?z?�?�?�/�/�. �:�?�;O??�?ZO lO~O�O�O�O�?�?�? �?O_5_(O:O�Oz_ �_�_�_�_�_�O�O�O� _"_4o `� @Ȁme�/{oW__Y�a�UDo�o�o�_�j �o�o1CaI� �gq����� ��Q�c���7�i��� ��������Տ�ُ�\�
�ol��A��*SYSTEM*��V9.10185� ��12/11/�2019 A ��� ��r�ӓSR�_T   � �$ĐENB_T�YP   �$RUNNER_�AXS� $HA�ND_LNGTH��`�THICK���FLIPґ�`�$INTFERE�NCE��IF_�CH��I֑$��9�INDXD�ĐG�1POS  � W�N�`�ANG�`�x�_JF��P�RM`� 	�R�V_DATAƑ�  $��ET�IME  ��$V�ALU����GR�P_   ���A  2 ��SCő	�� �$ITP_��� $NUM�ڠOUِ	�TOT��
�DSP!�JO�GLIM� $F�INE_PCNT�@�CO��$M{AX�TASK@��KEPT_MIR|=�]�PREMTq��}�APLD���_EX������t�@���PG��BRKHO�LD�!��I_��  ڲ@���P_�MADE�w�BS{OC�MOTN��DUMMY163��SV_CODE�_OPM�SFSP�D_OVRD��fR�LDL�O�ORZ�[TPӐLE[�F!�l[�:�OV=�SF�ʈᐓ�T�F��A�a�U�FRA��TOOL~@�LCHDLYW�RECOVK��:��WSs�:��=�RO�M��I�_�ڐ �@��S��NVER]T�OFS;�CǠD�FWDt���p���ENAB��7�TR���`���E_FD}O��MB_CM�z��B-�BL_Mi��]��Ҫ�2S�VST=AA�$UP���2��G�׸�AM����0а��%� �_M��A��AM�A�1�T$C�A0�,�D�7�HcBK���L�IO?��[�IQ�$PPAO�{�`��s��s�~1�DVC_DB�� F����쑼��A���1��%���3��+�ATIO� �h�K�aU��/�/�P�ABF�T֒E�G�Ԛ���E��:�_AUX�SU�BCPU�G�SICN_7Ў���P�1�������FLA��ݑHW_C1���j������$ATR���_$UNIT���>��ATTRI����G�CYCLC�NE�CA!�FLTR�_2_FIR�TARTUP_CN`�޶�SIGNO�LPxS�2�1�_SCTz�F_��F_��t���FSF����CHA���[���O��RS�D/���/�P��s�_T��PRO�|�p�GEMP�=��T�ę�ܐ���'DI�AG�RAILAiC��p�M�LO�4�'�4�PS-�@�� i�+�%�PR��S^B�  �C��� 	$�FUN�C���RINS�_TB���=�o�RA��`�7��a��E��WARq�8�BOLCUR�$A+	((DA��G(#%LD=�?�h�o#d��to#TI���%�ܐ$CE_�RIA_SWA�AF��P^��#��%�T2\CK��CM�OI���DF_L�E�_�PD�"LM���FA�HRDYYO��E�RGt H� �z���O 5MULS�E� ���0��$�JW�Jrǂ�FAN_ALMLV���1WRN�5HARDאO�_O,� ��2�1STO�Ƶ_,���AU��R�(���_SBR���5.��J���CMPINFڐ��-De!8C7REG@�NV0l�|$�۱DAL_N��sFL����$M �2��7%�ܐ�8�EC�M-�N0�Y���h��G���SP$R�W$Y��Z����|ۡ��� ����EG!`
�?�
QAR�0�'�20�U3 ��wAXE$�ROB!�7RED!�WR�߱_i]�SYܰDQ�:�VS�WWRI�V��STR �)��f�E��Ġ&To�1��B�P1��V5c�O�TOHAĠ�AR�Y�b]�ΡR�F�I��h�$LIN�K�!��3a$EXST_�S1�%U6�N[aXYZ�2ej7sf'OFF9�2bZbNh%`B���d�����cFI �g�hA�7Ĩ9�_JL��¢d�?ch��0�T�[8�US��B	qL2Ar�C7 ��DUO�$V9.pTUR�0X�#zu�!a(BX�P,�)wFL�[`��@�P�p|e�Y3y0�G� 1Ġ%KF�M�'�3��sp�����a�ORQ .���x��s��m�� ��H��,�_A]�OV	Ed���Mh l��C~� �C~��B}��0{�B�|� ��{�~��h� ��e� u�����l�v�e����0�C���.�ERK���	tEЪ��E�A�ܐ�e� gN!K�N!AX�¢N!� ��4b��0��Z1��o ��`��r`���`��:p��qp��1�p��:0�� :0��:0Ǚ:0י:0� :0��:0�:0�:0'��D�8�DEBU���$��3(�N�VbA!BNL�t�^�VA�� 
����+��� 7�0�7�o7�a7�ra 7��a7�:q7�qq�$Fp��"ۂ�cLAB�b8)�����GRO: )r�<*�B_,��T m��`�0��*���1�AND�pt�:�+�_e=��1Y� *��A�P`m�!|�- ^`NT�0ӟ�VELل���L���SERVE����@ $�`�A6]!��PO@ҹ ���`���@���!�@�  $�T�RQ�r
 �tR
����"2�q I_ 	 l���['ERR�boI,���لr�TOQلրL�HP���R�� G��%lHa��   �REP  
 ,��#�=��݁RA�� 2	 d��s��@���7 �@$r��� ����OC?!��  d�COU�NT�Q��FZN_wCFG	� 4��aF3T������ܣq �����AT��C �(�M��g2��Ճ{����FA� 䅻&��XdP�����SQ���G�dQPB����SHEL}@Y�� 5pB_B;AS��RSR`F�E^SS��!M�1�תM�2p�3p�4p�5*p�6p�7p�8��@�ROO�p��V ]`NL�ALsAB��FN�ACK�IN�T�g �CU�0E0� 	_cPUdq�2ZOU��P�aH-�֨ �P���TPFWD_KA1Rw�iAf�RE��$0qP/`U!w�QUE`I@ e�Up�r�0�1I�0��-�[`S��SF[aSCEM3��A�0A��7STYSO� 	�DI�}����!�_TMuCMANR�QL[`END�t�$KEYSWIT�CH^s.�HE�UpBEATM�PEPLEv������UrF�sS3D_O_HOM� O�16 EFA�PR�a�(vQ�P�EC�O01c���OV_Mr� � �IOCMGt�A��	P,�HK�A DHXabG��U^ҹMPx�W�WsFORCfC7WAR 2��@.��OMP  @���c�0U�SP3P1(�&�@�$3�&4���*�O� L�"��aHOUNLO9 \�4�ED�1  �S�NPX_ASZ�; 0�@ADD���$SIZfA$�VA���MULTKIP��.3� A�! � $H	�/0��`BRS}�ϱC<rТ6FRIFu��aS� �)��0NFOODBU�P~��5�30�9�ƽAfIA�!$V��y�x�R�SN��@� � L0��TE��s8�:sSGLZATAb�p&o�sC᳍P[@OSTMT�q�CPP�VBWe�\DSHO�W�Ev�BAN�@TP�`�wqs8��s8��r���V7�_G�� :p$PCD �7���kFB�!PXSP� �A U�ADP���� �W�A00^�ZR� bW� bW� �bW� bW5`Y6`Y7�`Y8`Y9`YA`YB�`Y� bW��cV�@bWF `X7�$hlY(@$h�Y@@T$h�Y1�Y1�Y1�YU1�Y1�Y1�Y1�YU1i1i1"i2_YU2lY2yY2�Y2�YU2�Y2�Y2�Y2�YU2�Y2�Y2�Y2�YU2i2i2"i3_Y��p�xyY3�Y3�Y3��Y3�Y3�Y3�Y3��Y3�Y3�Y3�Y3�i3i3"i4_Y4�lY4yY4�Y4�Y4��Y4�Y4�Y4�Y4��Y4�Y4�Y4�Y4�i4i4"i5_Y5�lY5yY5�Y5�Y5��Y5�Y5�Y5�Y5��Y5�Y5�Y5�Y5�i5i5"i6_Y6�lY6yY6�Y6�Y6��Y6�Y6�Y6�Y6��Y6�Y6�Y6�Y6�i6i6"i7_Y7�lY7yY7�Y7�Y7��Y7�Y7�Y7�Y7��Y7�Y7�Y7�Y7�i7i7"d��@Pz�U� ��߰e�
�A�2�� �x #�R�@  ��M��R9� ��Q_+�R����(�~ J��S/�C�D�^��_U�0i��"YSL|���� � L5 Bj��4A7�D����&RVALUj�% x�1���F��ID_L��3��HI��I�"$FILE_L!�i�$���SA�� h	�M�E_B�LCK�Z�uAc�D_CPUs�M0s�A0�u�$�6�-0YZ@FR�  � PaW-����0��LA�A�S�������RUN_FLG���� ���v�!���!���H`F ��C���CAT2x�_LI�"  ]��G_O�� �P_EDI�"�@T2��c�k�9��pnє0�0��BC2LT �Q@ �(0��!c�FT���	T�DC�A4z���M0�������TH�0�!�#�$�R��0e ERVE�F�	F��5A�� �  �X -$q�LE�N�~�	q�) RA�� 2��W_?���14q��2��MOk�5	S�0 I. Z������q���DE�1LgACE,":�CC3Z¶_MA20>>TCVEfTXg
�|
8RQ��QJAUMD���J>JP�
}�2��@BP	l0JKVK�A .)A.5A#J�AF�2JJ:JJBAAL2h:hbAA2f5#� N1��(XB G�L��_�AA��ٱm�CF62! `	�GROU��vA�2�$QN��C�3�RE�QUIR1��0EBqU�3m��$T 2 *!n�&��50���" \� ��APPmR  CLG�
$t��Ng(CLO��w)S���)
��u6# ���M �C � 2�$'_MGA� CLPN�p�(� R �'BRK�)�NOLD�&�@RTCMOb�:
=�%Jb�4Pj  :  B  P�  �  6W57W5�hA���$� "���A�7)A�3PATH�7�1�3�1����3� / #\�PS�CA�� 7h"�!INFp�UC����0@C:PKUM9HY��?��  @A��L�[J�0[Jq0[@�PAYLOA7J{2L�R_AN���CL�ЦI�A�I�A�%�R_F2LSHR@��ALO�D~A�G=C|�G=CACRL_�� -E P)G�D�H��G��$H�"NRFLE�Xj#k�J��% PT"����E�W�A�kP>p�& :}���  �W�T��� ������F1�QEeYg���� ��(�bE2D Vhz����`x }t��m`�x��H�QT�w^qXF� ��d�h%.�x1 CUgktb��С���J�' ������	/���A1Trf!� EL�`���D�#(J/ &* JE�0CTR)AmaTN���@�'HAND_�VBG�jQ���4(� $�pF2�&�f��SW���TB�&)� $$M�@ �)!��!�1�#p��E2�A���@�&��<���-A�,���*A;A�;G��+���*D;D�;P�0G��ݩST��'�9�N8DY �e �&(�O��@r��G �Q�G�A�G�t`�5P_5h5q5z5�5�5�5�3 �R�4* ��T�2 �a㵙!��ASYMEeP� F)K� L�A$O_ B�X5@HD2=4ĸ�ROdOvO�O�CJ�LR0�Jp�����Id_VI���ؙ#!�V_UN ���6�W��AJN� |�N��LR�U_ԃ�]�� $YR03_E_���d[TcS α��HR�����+���}P]"D�I0#O#���9���, g�V�I9�AV1SP�s`^��^�v`��ϰ�`� �- � ɑMEB�a��y���`�T�PT��Հ�0����AV �������T���� $DUM�MY1q1$PS�_p`RF2`��$����PFLA�Y�P���$GLB_T��1���]!�S��aq�}�. XXT '�1ST�* �SBR�0M21_�V&"T$SV_E�R�@O��w��CL�K�w�A�`OS� �G�L�EW�/ 4\���$Y��Z��!W���AœAz�9B�Υ0��U��0 ��pN���$G�I��}$�� �/�����1 qL���}$F�½ENEAR�`N�wcFd	�`TANC�wbͱJOG&`H0 �2Ӑ$JOI�NT�"��ҽ�MS�ET�3  EJ�a�S�����_4� n`U�a�?�* LOCK_�FO�@Б�BGL�Vt�GLTES�T_XMj �EM�P� &"2I�� c$U�P��9`20* ���X1#̐� X/�y�CE�&y $�KAR$qM%�TP�DRA���VE�C`�� IUX2�]HE TOOL�9c�V8dRE�I�S3�U�6z1m`ASCH� / 3�O@ԩ���3g�% SI�Z"  @$RAIL_BOXE����ROBO)?����HOWWAR�VQH!��!ROLM �n%ԁ$"�6 a`n�0O_F�!��HTML5�)AH��!�15�5�R�O�R6�1`�� ґv��OU�7 d���T/`�J�$�� $PIP*N�p�6"�!`X� �PCOR�DED� 
@� a XIT*0) � �O`� 8 D 0�OB|�N�� �7v1��p/�v2��P�SYSv1�ADRO� ��TC}H� 9 ,�pSEN	�QA_��4݁0���VWV�A|�: � �����PREV_�RT��$EDI}T(FVSHWR��c�G@�b���D��O�^DW�$H�EAD����x@���0CKE����CPS�PD�FJMP�0Ld�ϰR�`;�;~0T{Q�6I3SO�C���NE�P���TIC�K9c��M�QͲ�CH=NY�< @�0�AᅗA_GP&V-&�PgSTY�2!LOK����B"R�P= tk 
#@G�5%$A�=c�SE�!$@D�9`���M��P&�&VSQU�,e�яTERC����אS�>  o�� �p��q�``O����F{`IZ����PR\0�Db�A0P9U;�Te_DOi�0�XS� K�AXI4s`�#]UR��c@P�O P�6���_��2ET�bP�0	ŐԐ� 
�sPA�����9'[) ��S=R��?l�P� !���/u�Ay�/u*� /s8�/sH�uuj�uuz� uu���u�}���u�|���yC
��}C�}�ϕϸ�Ϲ�5�SSC3� o@ h��DS4P�/���SPJࡅAT�x� �UaP�B��A_DDRES�B3@�SHIF�O_2+CHO��1IR����TUR�I�� }A�CUSTO�d*��V�I>�B�2���8c�
2
 BV81da~�C \a�8A�rPC�a�P��C���b�bR�6���T�XSCREEx2Dz��QTINA��# Ӕ�A�a��ٰE T�A��8b�1��n� ��a�2�b�/@RROS�~ �0�@�o�v� UE�DF ����1
�S��1RSMPwgUe0�P抡�S_��=Ú���ȧ�=õaC���� [2EΐUEմGD⸢��D`GMT��L�p��a~�O�� B�BL_ W��~�HS �rPJ�O��V��LE�a�N �`�RwIGHj�BRD���ہCKGR����T�f0����WIDTH@#T@�b)!��i�MI� EY��}�I
2б m VR6 @aBACCKTQ�Ũ���sFOS1�LAB_q�?(��I �$�URT!E�"�ް��H>@� J 8��~ !_wA�h�R��� s(����U�O�~�%KP����Uv���9Ry!LUM�ØfNՀERV!1R�Ph j�L���`GEI�0O�`l2�@LP��b	E�Pf�)%�v�3؆��3�  2�50�60�70�8��R��?`h ����� !�S�PK�ݱUSR��M �<a���U(�F�O�PRI�amx  ���TRIP2!m�UNDO;�N �P �ye`!xepS�P�`�P Oc�\��CaG PT� �T��^�OS��s�R �`F�J��Z�P���� ����6Th�PU�Z�Q���ã�5UJ�OSFF([�R_���=O)� 1P���Z;�Q��GU�1P:��V�Q�`��SUB86R���SRT��taSR}� #cOR N��RAU(p��T����7��_&@�DT |�1p�8OWNM��4�$SRCQ�Ҡ�PDx(&rMPFIMTl��`ESPPab� ���eA�������A@n
�U `��WO[pr�4a�PCOP��$�`O�_- ��,1�WA3@CF� � Z��"�@l"+�� V�SHAD�OW�`��_UN�SCA��ʴD�GD!�1EGAC<�8�K�VCWp`>
�W� ,"w16�S$NER�cȷQ#+�C0cDRkIV6f�a_V/P��@m D��MY_UBY��kyV��UR��P�eA�� "�P_MT"LZkB�M]�$�@DEY��3EX7�^��MUb�@X]�V$��US���`�_R�����
��R���G�pPACIN�A�PRG�$�"��"��"ң�RE}�遚�c�H�"@�X �� G�P���� @�IR��@Y ��?�ӱ��	�qa�REb#SW� _A$�!�`W#B`O��ہQA�^3/rE��UePd�d��JHKjRZ��v:�P&q[0%��3EAP�7� j�^5��IMRCV
�[� ��OvPMj�C·�	�2��#�2REF6�F�6�1M0���c 50���:FAJFAKhE�6�?_ �:�H�;�pS��N'�a����I�\ �GR�ӵ`4�м�POU4W�"<Vk W 5U��2��$Ԑ��C`,��Y��U�2Q{�ՀUL6j�Z_ CO~��3[H EPNTZ�T���U���V�ђSQPL���U#�U���W����VIA_���]� ��`HD�����$JO��6��?$Z_UPL�W�Z|pW!e�QPSp�0��_LI��$EP EQ��k�a�QǑ΁���΀G\m�^� �0���aw� ��CACHLO:A�d�a�I �i��� 1CI`M%I�FHa�eT�p�fN�K$HOj��`OCOMM���Ot� wWӲ�S&�T7 �VP�"@�mr_SI	ZwtZ� rx!asw���MP�zFAIj!`G�4�`AD�y��MRET�r|wG�P��> & �ASY�NBUF�VRTaD�%�|q��OL��D_��A�W��PC&��TU7#�`Q{0	��ECCU�(VEM�� �e���gVIRC��q9�!���%�_DE�LA�#&Q���AuG5�RK!XYZ̠��K!W1��8A���2��TN8"IM߁8�������eGRABBJ��Yb" �e�_e��LAS��A�a_GE�e`u�&��;���T/S&N` ����%I���"ņ�BG2f�V5��PK� ǆ,�aWGI��N#�`2A�A@��`�qq�a+ⒹaS�p�fN:�]�LEX��b�����;��Nq��I? �-|�� |�.$�3k��- 
�"c��b�t�Ŀ�\�a�ORD����Qp��w�RN�d $MPTIT� �C���F�VSF����e�  -�[�QK URl�3]�SM!�f+���ADJ�N%�PZ�D>�g DƨBaA�L+`�p�AbPER�Is`��MSG_Q9�$}q�u���b��h+�"�g�J`�3p/�XVR#�in�b��T_OVRi���/ZABC��j�";�,s/@
 i�Z]�#�k+�=$L�-B��ZMPCF��l�H���A����LN�Kc�
^�MK!��m $,q�0�įCMCM� C�C����DP_A+A'$J����Dbq� ��� �� ����
D��F�UX���UXE]!f��	�]��]��oс�oё���FTF�sQӾ�A9�b�nC {�}����YJ`]D�� oY�R�p�U�$HEIGH�#"�?(MP�.A�����Dp � EX�$BQPx ��SHIF�s��R�VI`F��/B|�0�C `�dTF {"���蕓��WuD��TRA�CE��V�A^� P�HER� q �,MP�)�;��$�R�!p�� ����F��\� 6�S�F��  S�x�2p������s���r������	��U�C�AD�C��8l6�R  d�� ZD �Qx0C����l�l0�V| �6�V���@ 2F���� D� P����� 	�	F�,:$ZH ~l������ � //D/2/h/V/x/ �/�/�/�/�/�/
?�/ ??.?d?R?�?v?�? �?�?�?�?O�?*OO NO<OrO`O�O�O�O�O �O�O�O__8_&_H_ n_\_�_�_�_�_�_�_ �_�_�_4o"oXoFo|o jo�o�o�o�o�o�oF���$SAF_DO_PULSC�G��@k�$qp���|k����5qR ���`�X^P�\�\�[������s��[� ����� ���*�<�N�`�r�섏���  "��2��[���d��ȁq�rs�� @��@����*�܉�� � �6��_ @J�TY J���������?T D����� ���)�;�M�_�q� ��������˯ݯ��x~������M�_�$��sR�;�4�f���p����
�t��Di���q��  � � ���R�q|ulq�� �%�7�I�[�m�ϑ� �ϵ����������!� 3�E�W�i�{ߍߟ߱� ����������/�A� S�e�w�����S��G�������0�B� T�f�x�������� ������"4FK��b0E�ҳD�ܽ� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? ��?�?�?�?�?�?�? 	OO-O��QOcOuO�O �O�O�O�O�OLz� �!_3_E_W_i_{_�_ �_�_�_�_�_�Yoo ,o>oPoboto�o�o�o �o�o�o�o(: L^p�������ø��Ǔ�6� H�Z�l�~�������Ə ؏���� �2�D�V��d�#�m�����������i�	12345678ݲ�h!B!�)�Tz1!���
� �.�@�R�d�v����� ��"�ïկ����� /�A�S�e�w������� ��ѿ������)�;� M�_�qσϕϧϹ��� ������%�7���� m�ߑߣߵ������� ���!�3�E�W�i�{� ��L߱���������� �/�A�S�e�w����� ����������+ =Oas���� ���'9�� ]o������ ��/#/5/G/Y/k/ }/�/N�/�/�/�/�/ ??1?C?U?g?y?�? �?�?�?�?�?�/	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_"BS��]_o_�?�_��_�_ԚCz  �Bp�z   ���2�� } ��X
g�  	��R2U_<oNo`oro�l��\�+o�o�o �o�o"4FXj |������� ���oB�T�f�x��� ������ҏ����� ,�>�P�b�t�����������Qa�R<Ք� ˕a  �������#a#at  �P#�;����`�$SCR_�GRP 1��*P�3� �� ��R ��U	 ����������Qԑ �U������ٯǯ ��]g�`��C�,�����m��C����l�LR Mate� 200iD 5�67890!`L�RM|� 	LR�2D ���
1'234��Ц�d��hbճ���}�ݣ}��cԑ����ѡ�	j4�F�X�j�|τ�?��H������}���į������̦<��1��A���e���WV��Vh`,R���  W��B���Pư߮��Ԫ�A�P��  @�0�ժ�3@����� ?4��ª�H�P'��ڪ�F@ F�`Q�Y�P� }�h���������� ���ʩ�����J�5�G�Y�k�B�y���� ��������=( aL�p��o�
'�����W`�.�4�@4�>�7�4̧@��n�PQ�����ݣT_��AA�������aĲ�1 
/1/C/�Q*!f(r/�/S/�P�#
b�/�/�/�� ?�/$?,4]�ECL�VL  �1�����>1L_DE�FAULTF4���_��0Z3?HOTSTRf=��z2MIPOWER�FE0�Ur5�4W7FDOg6 r5=2�RVENT 1�M1M1�3 L!DUM_EIP,?�H�j!AF_�INEf0+O3D!�FTOZN!O~O!��ϣO �mO�O!�RPC_MAI�N�O�H��O_�CV�IS�O�I�_b_!7TPUPPUY_I�dQ_�_!
PMON_PROXY�_�Fe�_�_uR�_Mf��_Fo!RDM_'SRVGoIg5o�oG!R���oHh�o��o!
�@MoLi��o*!RLSY3NC+Qy8v�!ROS O�|�y4e�!
CEwP�MTCOM�Fk��!	�rCON�S�Gl�Z�!>�rWASRCaoF�mI���!�rUS	B��Hn���O� Uc���?�d�+���O��s�П87RVICE_KL ?%�;� (%SVC�PRG1ן�	�2��$��3G�L��4�o�t��5�����6��į�7�����$/�*�97�<���o d������9���� a�ܿ�������,� �ٯT���|��)� ���Q���6�z���6� ���6�ʿD�6��l� 6�ϔ�6�Bϼ�6�j� ��6����6���4�6� ��\�^�
�ܟ���� �����.������8� #�\�G���k������� ��������"F1 X|g����� �	B-fQ �u�����/ �,//P/;/t/�/q/ �/�/�/�/�/�/??�(?L?7?p?�_DE�V �9��UT1:|?�0GR�P 2
�5����bx 	� 
 ,�0x?�?�2�? OO@O'O9OvO]O�O �O�O�O�O�O�O_*_ _N_5_r_�_�?�___ �_�_�_o�_&o8oo \oCo�ogoyo�o�o�o �o�o�o4�_)j !�u����� ���B�)�f�x�_� ������������M� ,��P�7�t�[�m��� ��Ο�����(�� L�^�E���i������ ܯ�� ����6��Z� l�S���w�������� ѿ���2�D�+�hϿ� ]Ϟ�U��ϩ������� ��@�R�9�v�]ߚ� �ߓ��߷�������*� ��N�`�G��k��� ���������&�8�� \�C�����y������� ��C���4F-j Q������� �B)fx_ ��������/ ,//P/7/t/�/m/�/ �/�/�/�/?�/(??�!?^?e3d �e6	 L?�?�?�?�?�?�?O�K%�O5O<C���NA�1NE^OlGVO �OzO�O�O�O�I"O_ JI�O4_"_X_F_h_j_ |_�_�O�__�_o�_ 0ooToBodo�_�_�o �_�o�o�o�o, P�ow�o@�<� ����(�jO�� ���p�������܏ʏ  �B�'�f���Z�H�~� l�������؟���>� ȟ2� �V�D�z�h��� ��ůׯ��������.� �R�@�v�����ܯf� п������*��N� ��uϴ�>Ϩϖ��Ϻ� ������&�h�Mߌ�� ��nߤߒ��߶���.� T�%�d���X�F�|�j� ��������*��� ��.�T�B�x�f����� ���������* P>t�����d� ���&L� s�<����� �/T9/K//$/� l/�/�/�/�/�/,/? P/�/D?2?T?V?h?�? �?�??�?(?�?O
O @O.OPOROdO�O�?�O  O�O�O�O__<_*_ L_�O�O�_�Or_�_�_ �_�_oo8oz__o�_ (o�o$o�o�o�o�o�o Ro7vo jX� |����*�N �B�0�f�T���x��� ����&�����>� ,�b�P���ȏ����v� ��r�����:�(�^� ����ğN�����ȯʯ ܯ� �6�x�]���&� ��~�����Ŀƿؿ� P�5�t���h�Vό�z� �Ϟ����<��L��� @�.�d�R߈�v߬��� ��ߜ����<�*� `�N���߫���t��� ������8�&�\��� ����L����������� ��4v�[��$� |�����<! 3��T�x� ���8�,// </>/P/�/t/�/��/ /�/?�/(??8?:? L?�?�/�?�/r?�?�?  O�?$OO4O�?�?�O �?ZO�O�O�O�O�O�O  _bOG_�O_z__�_ �_�_�_�_�_:_o^_ �_Ro@ovodo�o�o�o �oo�o6o�o*N <r`���o� ���&��J�8�n� �����^���Z�ȏ�� �"��F���m���6� ��������ğ���� `�E����x�f����� ��������8��\�� P�>�t�b��������� $���4�ο(��L�:� p�^ϔ�ֿ�������� ����$��H�6�l߮� ����\��ߴ�������  ��D��k��4�� ������������^� C����v�d������� ����$�	������ <r`������  �$&8n \������� /� /"/4/j/��/ �Z/�/�/�/�/?�/ ?r/�/i?�/B?�?�? �?�?�?�?OJ?/On? �?bO�?rO�O�O�O�O �O"O_FO�O:_(_^_ L_n_�_�_�_�O�__ �_o o6o$oZoHojo �o�_�o�_�o�o�o �o2 V�o}�F hB���
��.� pU�����v����� ���Џ�H�-�l��� `�N���r�������ޟ  ��D�Ο8�&�\�J� ��n�����ݯ��� ���4�"�X�F�|��� ���l�ֿh����� 0��Tϖ�{Ϻ�DϮ� �����������,�n� Sߒ�߆�tߪߘ��� �����F�+�j���^� L��p�������� ������$�Z�H�~� l��������������  VDz��� ��j����
 R�y�B�� ����/Z�Q/ �*/�/r/�/�/�/�/ �/2/?V/�/J?�/Z? �?n?�?�?�?
?�?.? �?"OOFO4OVO|OjO �O�?�OO�O�O�O_ _B_0_R_x_�O�_�O h_�_�_�_�_oo>o �_eowo.oPo*o�o�o �o�o�oXo=|o p^������ 0�T�H�6�l�Z� |�~���Ə��,���  ��D�2�h�V�x�Ώ �ş�������
� @�.�d�����ʟT��� P�ί�����<�~� c���,���������ʿ �޿�V�;�z��n� \ϒπ϶Ϥ�����.� �R���F�4�j�Xߎ� |߲������ߢ��ߞ� �B�0�f�T���߱� ��z����������>� ,�b������R����� ��������:|�a ��*������ �Bh9xlZ �~����> �2/�B/h/V/�/z/ �/��//�/
?�/.? ?>?d?R?�?�/�?�/ x?�?�?O�?*OO:O `O�?�O�?PO�O�O�O �O_�O&_hOM____ 8__�_�_�_�_�_�_�@_%od_nQ�$SE�RV_MAIL � nUd`�JhO�UTPUTYh�oP@NdRV� 2�V  g`� (�Q4o�oNdSA�VEzlhiTOP1�0 2�i d j_ 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ����U�e�YP�oKcFZN_�CFG �U�gc�d�a�eT�G�RP 2^��a ,B   A��~nQD;� B����  B4�c�RB21�fHELLW��U�f�`�o�u���%RSR��)�b�M���q� ����ο��˿��(���L�7�pςϔ��/  �a%����P�Ϣ�����oP��L������Ǫ�2oP�d����ɦHK 1׫ ߈߃� �ߧ����������� %�7�`�[�m���������ìOMM �ׯ�ȢFTOV�_ENBYd�a�iH�OW_REG_U�I7�LbIMIOFWDL����l�/WAIT4���v�Ȕ�t`X��d��TI�MX�����VA�X`��l�_UNIT�3��iLCQ�TR�YX��eN`MO�N_ALIAS k?e��`heo �����
t�� #�GYk}� :������/ 1/C/U/g//�/�/�/ �/l/�/�/	??-?�/ Q?c?u?�?�?D?�?�? �?�?O�?)O;OMO_O qOO�O�O�O�OvO�O __%_7_�O[_m__ �_�_N_�_�_�_�_o �_3oEoWoioozo�o �o�o�o�o�o/ A�oew���X ������=�O� a�s��������͏ߏ ����'�9�K���o� ��������b�۟��� ���"�G�Y�k�}�(� ����ůׯ鯔��� 1�C�U� �y������� ��l����	��ƿ?� Q�c�uχ�2ϫϽ��� ���Ϟ��)�;�M�_� 
߃ߕߧ߹�d����� ��%���I�[�m�� ��<����������� !�3�E�W�i������ ����n�����/���Sew�����$SMON_DE�FPROG &������ &*SYS�TEM*�� �	�RECALL� ?}�	 ( ��}xyzra�te 61=>192.168./�07:15032} . 36 2T�Zl~�}
!11 ,>P��/ � ���g/y/�/� }9copy �frs:orde�rfil.dat� virt:\tmpback\+/�=!�/�/�/�0�"m?db:*.*�/�/A �/c?u?�?�5�/�(emp;>254�4 W?�?�?O}-�6*.d�?�>�?aO8sO�O�61 ,O>O PO�O�O_�!/�:@�O�Oc_u_�_�1!4�:prog_1.tp�O�<S_�_�_o�8�?�/�_�PYoko}o�M/!?<o4ZRo�o��o�3x!d:\ �o+p�o�P�ofx�
�4!ua);�Y� ��o"o4o��i� {���o;��oV������ }6!��??;1052 ؏i�{��.!O;�M�P���� �O�O��Ο_�q���/ (_Q�A�S������/ -���N�Z�l�~�?�� >�M�R����Ϛt!��3�?41.15:8892Ѐؿi�{��,��;�M�O������ �)�����^�p߂����J�?�Q��������tpdisc 0��2 ����`��r���tpconn 0�3�E�W� �����������a�ps������Qick�_�=�P�������drop������bt� ��<?&FX��� ����gy�� 0BT��	/� ��c/u/�/�,/>/ P/�/�/?/*/�/�/ _?q?�?�/�/:?L?�?�?O�7!�3��?;� ZOlO~O��>O��RO��O�O_��$SN�PX_ASG 2����,Q�� P 0 �'%R[1c]@L�_WY?��%W_�_f_�_�_�_�_ �_�_o�_7oo,omo Powo�o�o�o�o�o�o �o3W:L� p�������  �'�S�6�w�Z�l��� �����Ə����=�  �G�s�V���z���͟ ��ן��'�
��]� @�g���v�������� Я��#��G�*�<�}� `�������׿��̿� ��C�&�g�J�\ϝ� �ϧ��϶�������-� �7�c�F߇�j�|߽� ������������M� 0�W��f������ �������7��,�m� P�w������������� ��3W:L� p������  'S6wZl� ����/��=/  /G/s/V/�/z/�/�/ �/�/?�/'?
??]? @?g?�?v?�?�?�?�?��?�?#ODTPAR�AM ,U�6Q �	�'JP�'D�@'H~D��-PPOFT_K�B_CFG  �fC2USOPIN_�SIM  ,[�sF�O�O�Ov@=@RV�NORDY_DO�  }E�ERQSTP_DSB�N�sBU_aX=@SR ��I � &ȃE�_�\�T�CTO�P_ON_ERR�_;B�QPTN ��E�P�C��RRING_PR�M�_0RVCNT_�GP 2�E�A�@x 	Q_Poh@>o�wobo�olWVD%`ROP 1LI�@�a xI�g�o�o�oE BTfx���� �����,�>�P� b�t�������яΏ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�]�Z�l�~��� ����Ưد���#� � 2�D�V�h�z������� ¿����
��.�@� R�d�vψϯϬϾ��� ������*�<�N�u� r߄ߖߨߺ������� ��;�8�J�\�n�� ������������ "�4�F�X�j�|����� ����������0 BTf����� ���,SP�bt����bPRG_COUNT�Fs��R�ENBo��M��D/_UP�D 1{[T  
�gBR/d/v/�/ �/�/�/�/�/�/?/? *?<?N?w?r?�?�?�? �?�?�?OOO&OOO JO\OnO�O�O�O�O�O �O�O�O'_"_4_F_o_ j_|_�_�_�_�_�_�_ �_ooGoBoTofo�o �o�o�o�o�o�o�o ,>gbt�� �������?� :�L�^���������Ϗ ʏ܏���$�6�_� Z�l�~�������Ɵ������_INFO� 1@%& H�	 �c�N����r�?�2@B?�z=��t���"�DA�/�?������µ�B�QQ���=�@ @G� A�i��>�| >���� �D�b�����B��B�3�~ՠS�B�����²�B����j�r7菟5B��/��Y?SDEBUG�A ���d))Q�SP_�PASS�B?~c�LOG =�]J!  �����  �%!�UD1:\��#���_MPC��@%�#ϒ@!̱A� @!�SAV ���y�ظ�вC�׸SV��TEM_TIM�E 1��K � 0  ����C�CȀ�	��MEMBK  @%�%!����%�7�G�wX|& � @G���iߎߞ�b��߲����^� y�@ ����*�<�v�T�f�`x������ ��� ����
��.�@�R�d�v��e���������� ��(:L^p ������� ��SK�����@hRdX�� "�Q2sߣ�P� �� �������%/7/I/[/O�u$� �u/���@�/�/�/���/�À?@'?9?K?]?o?�$s?�?���?�4^�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__�)�T1SVGUNwSPDy� 'c���4P2MODE_?LIM ��g�20T2=P]Q��/U�ASK_OPTI�ONX��g��Q_�DIr�ENB  ���c��QBC2_?GRP 2#c�0���_�"� C�c(\�BCCFG !��[~� o"Ekem`eo���o�o�o�o �o�o�o?*c N`������ ���;�&�_�J��� n�����ˏݏ��ɋ�� ɏ*�<����r�]��� ����H�ڟԯ��� ��,��P�>�t�b��� ����ί������ :�(�J�p�^������� ��ܿʿ�� �6�� �J�\�zόϞ���� ���������.�@�� d�R߈�v߬ߚ߼߾� �����*��N�<�r� `����������� ��$�&�8�n�\��� HϪ���������|�" 2XF|��n ����� 0fT�x��� ��/�,//P/>/ t/b/�/�/�/�/�/�/ ��
??:?L?^?�/�? p?�?�?�?�?�? O�? $OOHO6OlOZO|O~O �O�O�O�O�O_�O2_  _B_h_V_�_z_�_�_ �_�_�_�_�_.ooRo ?jo|o�o�o�o<o�o �o�o<N`. �r������ �&��J�8�n�\��� ����ȏ���ڏ��� 4�"�D�F�X���|��� hoʟܟ������B� 0�R�x�f��������� �ү���,��<�>� P���t�����ο��� ��(��L�:�p�^� �ςϤϦϸ������ ȟ*�<�Z�l�~��Ϣ� �߲�������� ��� D�2�h�V��z��� ������
���.��R� @�b���v��������� ����N<r (ߊ����\��8&\Fz��$TBCSG_G�RP 2"F�  �z� 
 ?�   ��������@5//Y/k+~�$��d@ ��!?>z	 HBLk(z��&j$B$  C�`��/�(�/�/Cz�/�(=A�k(333?&ff?��i%�A��/m?80 k(c�͎6S5�0DHp?�=@�H0j%K1�5j$�1D"N!�?�?�?�? ;OJ�(I&�(nE�OLO ^O�O�O�O�O�O_ [��H:Q	V3.�00�	lr2d S	*\PTTy�k_*_ �Q�I 8�Pt]�_  �_�_,�[~J2�%�=Q�o�UCFG '�F� �"j��Lb�ROlwl�wo�o�jO�o�o�o �o�o=(aL ^������� ��9�$�]�H���l� ����ɏ��Ə���#� �G�Y��� d�v��� 2�����˟�ܟ� � 9�$�]�o�����N��� ��ۯƯ��zf6� BF�H�Z���~����� ؿƿ����2� �V� D�z�hϞόϮϰ��� �����
�@�.�d�R� tߚ߈߾߬����ߴ ����>�`�N��r� ����������&� ��6�8�J���n����� ����������"2 4F|j���� ���B0f T�x����� /�,//P/>/`/�/ 0�/�/�/l/�/�/? ??L?:?p?^?�?�? �?�?�?�?�?O O"O HOZOlO&O|O�O�O�O �O�O�O_�O_ _2_ h_V_�_z_�_�_�_�_ �_
o�_.ooRo@ovo do�o�o�o�o�o�o�o *�/BT� �������� 8�J�\��l������� ��ڏ����ʏ4�"� X�F�h���|�����֟ ğ���
���T�B� x�f���������Я�� ���>�,�b�P�r� t�����6Կ����� (��8�^�Lς�pϦ� �������� ߾�$�� H�6�X�~ߐߢ�\�n� �������� ��D�2� T�z�h�������� ������
�@�.�d�R� ��v����������� ��*N`
�x� �F���� $J8n��Pb ����/"/4/F/  /j/X/z/|/�/�/�/ �/�/?�/0??@?f? T?�?x?�?�?�?�?�? �?�?,OOPO>OtObO �O�O�O�O�O�Ol� _._�O_L_^_�_�_ �_�_�_�_ oo$o6o �_ZoHojolo~o�o�o �o�o�o�o2 V Dfhz���� ���
�,�R�@�v� d���������ΏЏ� ��<�*�`�N����� @_����ҟ|���&� �6�8�J���n����� ȯگ�����"��F��0�  l�p� �p���p��$TB�JOP_GRP �2(8���  ?�p�	�����*���@���@�� 0��  �� � � � ��p� @�l���	 �BL �  �Cр D�����<��E�A�S�<��B$�����@��?�33C�*���8œϞ�� �2�T�����;�2��t��@��?���zӌ�-�kA�>�Ⱥ�� �����l�>�~�a�s��;��pA�?��ff@&ff?�#ff�ϵ�8� ��L����}������:v,����?L~�}ѡ�D�H��5�;�M�@�33`�����>��|օ���8���`ự�	�D"��������`��r�|���"�9������g�v��x��� �������������� 0(V�b������p�C��p�	���	V3�.0�	lr2d��*b��k�p�{ E8� �EJ� E\� �En@ E��E��� E�� E��� E�� E��h E�H E��0 E� EϾ��� E���� E�x E��X F��D��  D�` E��P E�$��0�;�G�R��^p Ek�ui������(��� E�����?X 9�IR4! �H%�
z�`/r"�p�v#Ѭ߱/��E?STPARSI d�쵰��HR� ABL�E 1+��J p��(�' �k)�'��(�(o�w��'	��(
�(�(5p���(�(�(K!�#RDI�/��??(?:?L?^5�4O�?�;�? �?O O2N�"S�?�� �:�O__)_;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo���@ �O��7�isO�O�O�O U?g?y?�?�?�8�"pb�NUM  8�U����x� J �K �"_CFG �,Y{s�@��IM?EBF_TT�!u8��� �vVERI#�az�v�sR 1-�+O 8mp�k�2� ;��o  �� �,�>�P�b�t����� ����Ώ�����(� :���^�p��������� ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�{�V�h� ��������¿Կ���H
��"�q_Sq�v@�u�� MI_CHA�N�w �u u�DB'GLV���u�u�!�x�ETHERADW ?�%���v ��������(x�R�OUT�p!WJ!�*�H��SNMA�SK���s��255.��N�ߖߨ�N�� OOLOFS_�DI� BŪ�OR�QCTRL .�{>Cw/&�T�J�\� n����������� ���"�4�F�X�j�z���������#PE_�DETAI����P�GL_CONFI�G 4Yyiq���/cell/$�CID$/grp1��;M_q�9C�߮���� �,>Pbt� �����/�� :/L/^/p/�/�/#/�/ �/�/�/ ??�/6?H? Z?l?~?�??1?�?�? �?�?O O�n}�?VO hOzO�O�O�Oq���O�M��?__1_C_U_ g_�?�_�_�_�_�_�_ t_	oo-o?oQocouo o�o�o�o�o�o�o�o );M_q � �������%� 7�I�[�m������� Ǐُ�����!�3�E� W�i�{������ß՟ ������/�A�S�e� w��������ѯ������ �Us�er View �)	}}1234567890J�\�n����������5�	̿��0�2=���� �2�@D�V�h�ǿٿ7�3� �����������o�1�߾4��j�|ߎߠ߲���#���߾5Y��0�B�T�f�x��ߙ�߾6 ���������,���M�߾7��������� ����?�߾8u�: L^p������� lCamera;�1� 0BT2BE�~ ��H�����//�  ���f/ x/�/�/�/�/g�/�/ ?S/,?>?P?b?t?�?�����?�?�?�? OO,O�/PObOtO�? �O�O�O�O�O�O�?�7 XىO>_P_b_t_�_�_ ?O�_�_�_+_oo(o :oLo^o_�72+�_�o �o�o�o�o�_*< N�or����� so���a�(�:�L� ^�p��������܏ � ��$�6���7t� ͏��������ʟܟ��  ��$�o�H�Z�l�~� ����I��7(	9�� � �$�6�H��l�~��� ۯ��ƿؿ���ϵ�ǧ9��O�a�sυϗ� ��P������Ϙ��'�@9�K�]�o߁�
	�0߼��������� ��:�L�^�߂��� ������ߕ�� ��� 5�G�Y�k�}���6�� ����"���1C U���I+����� �����1C� gy����h�� �;X//1/C/U/g/ �/�/�/��/�/�/ 	??-?��![�/y? �?�?�?�?�?z/�?	O Of??OQOcOuO�O�O @?��k0O�O�O	__ -_?_�?c_u_�_�O�_ �_�_�_�_o�O��{ �_Qocouo�o�o�oR_ �o�o�o>o);Mx_qm  i ���������0�B�T�f�    v~������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ�ؿj�  
`( � �p( 	 ���B�0�f�T� ��xϚϜϮ���������,���� � �oq߃ߕ������� ����c`�=�O�a� �߅��������&� ��'�n�K�]�o��� ������������4� #5GYk����� ����1 C�gy���� ���	/P-/?/Q/ �u/�/�/�/�/�// (/??)?p/M?_?q? �?�?�?�/�?�?�?6? O%O7OIO[OmO�?�O �O�O�?�O�O�O_!_ 3_zO�Oi_{_�_�O�_ �_�_�_�_oR_/oAo So�_wo�o�o�o�o�o o�o`o=Oa s���o�o��� 8�'�9�K�]�o�� �������ۏ���� #�5�|�Y�k�}�ď�����şן���B�"�@� �*�<�N���$����+frh�:\tpgl\r�obots\lr�m200id��_�mate_��.xml
���Ưد����� �2�D�V�F��� `���������Ϳ߿� ��'�9�K�b�\ρ� �ϥϷ���������� #�5�G�^�X�}ߏߡ� ������������1� C�Z�T�y������ ������	��-�?�V� P�u������������� ��);R�Lq ������� %7NHm� ������/!/�3/E.g��� |$�r�<< p� ?�E+�/E/�/�/ �/�/�/?�/?<?"? 4?V?�?j?�?�?�?�?��?�?�?
O8OF���$TPGL_OUTPUT 7P��P� h  tE�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo�'otEh �=@2345678901Lo ^opo�o�o�o�cF�Io �o�o�o/�o3@ew���Ez}� ����'���]� o���������O�ŏ� ���#�5�͏C�k�}� ������K�]����� �1�C�۟Q�y����� ����Y�ϯ��	��-� ?�ׯ�u��������� Ͽg�ݿ��)�;�M� �[σϕϧϹ���c� u���%�7�I�[��� iߑߣߵ�����q��߀�!�3�E�W���HA} c!�������������@j/�.�p* ( 	 1oc�Q��� u��������������� )M;q_�� �����7 %GI[��?f�f &��-�#/ 5//Y/k/9j��/�/ H/�/�/�/�/?,?�/ 0?b?�/N?�?�?�?�? �?>?�?O�?OLO^O 8O�O�O�?|O�O�OvO  __�O_H_�O�O~_ �_*_�_�_�_�_�_o l_2oDo�_0ozoTofo �o�o o�o�o�o�o. @dv�o^�� X����*��� `�r����������ޏ <�N��&���2�\�6� H��������ڟt�Ɵ �"���F�X���@��� (�z�į֯�����j� ��B�T��x���d��� ���0���Ϣ��>� �*�tφ�俪ϼ�Vπ��������(�:��)�WGL1.XM�L��o��$TPOFF_LIM �|���}��N_SV��  �����P_MON7 8������2y�STRT?CHK 9�������VTCOM�PAT��6��VW�VAR :��\Y�� � q�������_DE�FPROG %���%MAIN� DT-��u�_D?ISPLAY�������INST_MSwK  �� ��?INUSER,����LCK5���QUI�CKMENY���S7CREx��7�?tpsc��5�Г���ҩ�_��ST�*��RACE_C_FG ;��Y�u��	z�
?���?HNL 2<��`� ��L^p�������
��IT�EM 2=8 ��%$12345�678901 � =<)Oai G !ow��3 �z��A//w )/��v/��/��/ �/M/=/O/a/{/�/�/ �/U?{?�?�/�??'? 9?�?]?	O/OAO�?MO �?�?�?qO�O#O�O�O YO_}O�OX_�Os_�O �_�__�_1_�_og_ 'o�_7o]ooo�_{o�_ 	oo�o?o�o#�o G�o�o�oSk� �;�_q:��U� �y�������%�� I�	�m��?�ŏ��Ǐ ُ���w�!�͟�� i�)�������+�՟�� �����ůA�S�e�� 7���[�m�ѯy���� п+��O��!υ�7� ������߿��ϯ��� ��K���oρϓ�߷� c߉ߛ��Ͽ�#�5�G� ����}�=�O��[��� �߲����1����g�����f���S��>|k��  ��k� ����
 ���������UoD1:\&��}��R_GRP 1?�� 	 @��q�m��������  ��&J5nY?�  ������� /�//'/]/K/�/�o/�/�/�/�/�/�/	�9�?%?{�SCBw 2@�� t q?�?�?�?�?�?�?�?�Oq�UTORIAL A��LOv��V_CONFIG B����	�O�[MOUTPUT �C���@�� �O�O__1_C_U_g_ y_�_�_�_�_�_�A�O �_oo1oCoUogoyo �o�o�o�o�o�_�o	 -?Qcu�� ����o���)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ� ���������'�9� K�]�o߁ߓߥ߷��� �������#�5�G�Y� k�}���������� �O�E�O'�9�K�]�o� ���������������� ��#5GYk}� ������ 1CUgy��� ����	/-/?/ Q/c/u/�/�/�/�/�/ �/�/?/)?;?M?_? q?�?�?�?�?�?�?�? O?%O7OIO[OmOO �O�O�O�O�O�O�O_  O3_E_W_i_{_�_�_ �_�_�_�_�_o_/o AoSoeowo�o�o�o�o �o�o�oo+=O as������ ���&9�K�]�o� ��������ɏۏ���|������0� B�,��m�������� ǟٟ����!�3�E� W�i��������ïկ �����/�A�S�e� w���������ѿ��� ��+�=�O�a�sτ� �ϩϻ��������� '�9�K�]�o߀ϓߥ� �����������#�5� G�Y�k�}�ߡ���� ��������1�C�U� g�y������������ ��	-?Qcu �������� );M_q�� �����//%/ 7/I/[/m//��/�/ �/�/�/�/?!?3?E?�W?i?{?�;�$TX�_SCREEN �1DD��,��}ipnl�/�0gen.htm�?�?�?OO%O���Panel �setup)L}��)OjO|O�O�O�O�O XONO�O__1_C_U_ �Oy_�O�_�_�_�_�_ �_n_�_-o?oQocouo �o�_,o"o�o�o�o )�oM�oq�� ���BT��%� 7�I�[�� ������ Ǐُ���t�!���E��W�i�{�������>U�ALRM_MSG� ?�9��0  ���*��5�(�Y�L� }�p�������ׯʯ�����ӕSEV  ��Q�ђEC�FG F�5�1  �%@� � A��   B��$
  ��#�5�� ƿؿ���� �2�D��V�h�v�]�GRP �2Gg� 0�&	� ����ӐI_B�BL_NOTE �Hg�T�G�l�"�0�!s�~��DEFPROݐ=%� (%�:� � (�a�L߅�pߩߔ� �߸������'��K����FKEYDAT�A 1I�9��p v��&�ϰ���0��������,(�+���$(POINT�  ]3�5���NC�EL_����NDI�RECT���� EXT STEP���6�TOUCHU����ORE INFOOaH �l�������9 ]o ���/frh/�gui/whit�ehome.pn�gp������}�point��*/</N/`/r/&  �FRH/FCGT�P/wzcancel/�/�/�/�/�/��#�indirec/4?F?X?j?|?�/� nex#?�?�?�?��? O$�touchup�?<ONO`O�rO�O$�arwrg�?�O�O�O�O_ �8#_5_G_Y_k_}_�_ _�_�_�_�_�_o�_ 1oCoUogoyo�oo�o �o�o�o�o	�o? Qcu��(�� �����;�M�_� q�������~��ӏ� ��	��-�4�Q�c�u� ������:�ϟ��� �)���;�_�q����� ����H�ݯ���%� 7�Ư[�m�������� D�ǿ����!�3�E� Կi�{ύϟϱ���R� ������/�A���S� w߉ߛ߭߿���`��� ��+�=�O���s�� ������\����� '�9�K�]��������з�����v���>����# 5WiC,U� M������ <N5rY��� ���/�&//J/ 1/n/�/g/�/�/�/�/ ���/?"?4?F?X?g� |?�?�?�?�?�?�?w? OO0OBOTOfO�?�O �O�O�O�O�OsO__ ,_>_P_b_t__�_�_ �_�_�_�_�_o(o:o Lo^opo�_�o�o�o�o �o�o �o$6HZ l~����� �� �2�D�V�h�z� �����ԏ���
� ��.�@�R�d�v���� ����П������/ <�N�`�r��������� ̯ޯ���&���J� \�n�������3�ȿڿ ����"ϱ�F�X�j� |ώϠϲ�A������� ��0߿�T�f�xߊ� �߮�=��������� ,�>���b�t���� ��K�������(�:� ��^�p����������� Y��� $6H�� l~����U��� 2DV-��X�-�������}���,�/
/�/.//R/d/ K/�/o/�/�/�/�/�/ ??�/<?#?`?r?Y? �?}?�?�?�?�?�?O �?8OJO)�nO�O�O�O �O�O��O�O_"_4_ F_X_�O|_�_�_�_�_ �_e_�_oo0oBoTo �_xo�o�o�o�o�o�o so,>Pb�o ������o� �(�:�L�^�p���� ����ʏ܏�}��$� 6�H�Z�l��������� Ɵ؟����� �2�D� V�h�z�	�����¯ԯ ������.�@�R�d� v���_O����п��� ��*�<�N�`�rτ� ��%Ϻ��������� ��8�J�\�n߀ߒ�!� �����������"�� F�X�j�|���/��� ����������B�T� f�x�������=����� ��,��Pbt ���9��� (:�^p�� ��G�� //$/ 6/�Z/l/~/�/�/�/��/���+�������/?=�/7?I?#6,5Oz?-O�? �?�?�?�?�?�?O.O ORO9OvO�OoO�O�O �O�O�O_�O*__N_ `_G_�_k_�_�_���_ �_oo&o8oG/\ono �o�o�o�o�oWo�o�o "4F�oj|� ���S���� 0�B�T��x������� ��ҏa�����,�>� P�ߏt���������Ο ��o���(�:�L�^� ퟂ�������ʯܯk�  ��$�6�H�Z�l��� ������ƿؿ�y��  �2�D�V�h����Ϟ� �����������_�.� @�R�d�v�}Ϛ߬߾� ��������*�<�N� `�r��������� �����&�8�J�\�n� ����!����������� ��4FXj|� ����� �BTfx��+ ����//�>/ P/b/t/�/�/�/9/�/ �/�/??(?�/L?^? p?�?�?�?5?�?�?�?� OO$O6O�8K}�����aO@sO�M]O�O�O�F,�_ �O�__�O2_D_+_h_ O_�_�_�_�_�_�_�_ �_oo@oRo9ovo]o �o�o�o�o�o�o�o *	�N`r��� �?�����&�8� �\�n���������E� ڏ����"�4�ÏX� j�|�������ğS�� ����0�B�џf�x� ��������O����� �,�>�P�߯t����� ����ο]����(� :�L�ۿpςϔϦϸ� ����k� ��$�6�H� Z���~ߐߢߴ����� g���� �2�D�V�h� ?������������ 
��.�@�R�d�v�� �������������� *<N`r�� �����&8 J\n���� ����"/4/F/X/ j/|/�//�/�/�/�/ �/?�/0?B?T?f?x? �??�?�?�?�?�?O O�?>OPObOtO�O�O 'O�O�O�O�O__�O :_L_^_p_�_�_�_}���[�}�����_�_�]�_o)of,Zo~oeo�o �o�o�o�o�o�o2 VhO�s�� ���
��.�@�'� d�K�����yﾏЏ� ���'_<�N�`�r� ������7�̟ޟ�� �&���J�\�n����� ��3�ȯگ����"� 4�ïX�j�|������� A�ֿ�����0Ͽ� T�f�xϊϜϮ���O� ������,�>���b� t߆ߘߪ߼�K����� ��(�:�L���p�� ������Y��� �� $�6�H���l�~����� ���������� 2 DV]�z���� ��u
.@R d������� q//*/</N/`/r/ /�/�/�/�/�/�// ?&?8?J?\?n?�/�? �?�?�?�?�?�?�?"O 4OFOXOjO|OO�O�O �O�O�O�O�O_0_B_ T_f_x_�__�_�_�_ �_�_o�_,o>oPobo to�oo�o�o�o�o�oh��{������ASe}=��sv,���}� ���$��H�/�l� ~�e�����Ə؏���� � �2��V�=�z�a� ������ԟ����
��� .�@�R�d�v����o�� ��Я�������<� N�`�r�����%���̿ ޿��ϣ�8�J�\� nπϒϤ�3������� ���"߱�F�X�j�|� �ߠ�/���������� �0��T�f�x��� ��=���������,� ��P�b�t��������� K�����(:�� ^p����G� � $6H�l ~������� / /2/D/V/�z/�/ �/�/�/�/c/�/
?? .?@?R?�/v?�?�?�? �?�?�?q?OO*O<O NO`O�?�O�O�O�O�O �OmO__&_8_J_\_ n_�O�_�_�_�_�_�_ {_o"o4oFoXojo�_ �o�o�o�o�o�o�o�o 0BTfx� �������,�@>�P�b�t���]����]������ÏՍ����	��, ��:��^�E�����{� ����ܟ�՟���6� H�/�l�S�������Ư ���ѯ� ��D�+� h�z�Y����¿Կ� ����.�@�R�d�v� ��ϬϾ�������� ��*�<�N�`�r߄�� �ߺ���������� 8�J�\�n���!�� �����������4�F� X�j�|�����/����� ������BTf x��+���� ,�Pbt� ��9���// (/�L/^/p/�/�/�/ �/���/�/ ??$?6? =/Z?l?~?�?�?�?�? U?�?�?O O2ODO�? hOzO�O�O�O�OQO�O �O
__._@_R_�Ov_ �_�_�_�_�___�_o o*o<oNo�_ro�o�o �o�o�o�omo& 8J\�o���� ��i��"�4�F� X�j��������ď֏ �w���0�B�T�f� ����������ҟ����� ���� ���!�3�E��g�y�S�,e���]�ί�� ���(��L�^�E� ��i�������ܿÿ � ���6��Z�A�~ϐ� wϴϛ������/� � 2�D�V�h�w��ߞ߰� �������߇��.�@� R�d�v������� ������*�<�N�`� r�������������� ��&8J\n� ������ �4FXj|� �����/�0/ B/T/f/x/�/�/+/�/ �/�/�/??�/>?P? b?t?�?�?'?�?�?�? �?OO(O��LO^OpO �O�O�O�?�O�O�O _ _$_6_�OZ_l_~_�_ �_�_C_�_�_�_o o 2o�_Vohozo�o�o�o �oQo�o�o
.@ �odv����M ����*�<�N�� r���������̏[��� ��&�8�J�ُn��� ������ȟڟi���� "�4�F�X��|����� ��į֯e�����0��B�T�f��$UI_�INUSER  �������  g��k�_MENHIS�T 1J���  (���?@(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1���+�=�Oπ9)��631Ϝ�������a�s�edi=t��MAIN�� �82�D�V� �'��v΁2ϡ߳������� ����%�7�I�[��� ��������h��� �!�3�E�W���h���@������������{� ۱{�*<N`r u������� &8J\n� �������"/ 4/F/X/j/|//�/�/ �/�/�/�/�/�/0?B? T?f?x?�??�?�?�? �?�?O��>OPObO tO�O�O�?�O�O�O�O __�O:_L_^_p_�_ �_�_5_�_�_�_ oo $o�_HoZolo~o�o�o 1o�o�o�o�o 2 �oVhz���? ���
��.�O+O d�v����������� ���*�<�ˏ`�r� ��������̟[��� �&�8�J�ٟn����� ����ȯW�����"� 4�F�X��|������� Ŀֿe�����0�B� T�?�Q��ϜϮ����� �����,�>�P�b� ��ߘߪ߼������� ���(�:�L�^�p��� ����������}�� $�6�H�Z�l�~���� ������������ 2�DVhze���$�UI_PANED�ATA 1L����� � 	�}/f�rh/gui�d�ev0.stm �M?connid�=0 height=100&_� �ice=TP&_�lines=15�&_column�s=4� font�=24&_page=whole� ��h�)prim/X  }[�0���� )�� �#/
/G/Y/@/}/d/ �/�/�/�/�/�/?�/�1?h��� �    ��in?�?�?�?�? �??�?_O"O4OFO XOjO�?�O�O�O�O�O �O�O�O__B_T_;_�x___�_�_�_�_E7  � �U�Oo$o6oHo Zolo�_�oO�o�o�o �o�ouo2D+h O������� 
���@�'�d�v��_ �_����Џ���Y� *��oN�`�r������� ��!�ޟş��&�8� �\�C�����y����� گ�ӯ�����F�X� j�|������ĿֿI� ����0�B�Tϻ�x� _ϜϮϕ��Ϲ���� ��,��P�b�I߆�m� ���/������(� :�L��p�㿔��� ������U��$��H� /�l�~�e��������� ������ DV�� �ߌ�����9 
}�.@Rdv� �����// �</#/`/r/Y/�/}/ �/�/�/�/cu&?8? J?\?n?�?�/�?�?) �?�?�?O"O4O�?XO ?O|O�OuO�O�O�O�O �O_�O0_B_)_f_M_�_�/?}��_�_�_�_
oo.o)�_So�5 Boo�o�o�o�o�o@o �o�o!W>{ b���������/��83;�$U�I_POSTYP�E  5?� 	 ;����a�QUICKME/N  p�����c�RESTORE� 1M5�  �*default�;�SINGLE~ԍPRIMԏ�mmenupage,23,1<� n�������G���П� ������<�N�`�r� ���"������ϯ�� 
��.�@��d�v��� ����O�п����� ï%�7�Iϻ��ϖϨ� ����o�����&�8� J���n߀ߒߤ߶�a� ������Y�"�4�F�X� j���������y� ����0�B�����a� s������������ ��,>Pbt�������SCR�E��?���u1sc�u2�!3!4!5!6�!7!8!�TATl�� ă5Y��USERTL#ks+�4�U5�6�7�8��a�NDO_CFG� Np��P�Qa�O�P_CRM5  ��U&a�PDd���Non�e���_INFOW 1O5f 0%��/�8o/�/�/ �/�/�/
??�/@?#? d?v?Y?�?�?�?�?���S!OFFSET Rp�j!�?��� �!O3OEOWO�O{O�O �O�O�OO�O___ J_A_S_�_w_�_�_�Kŏ�]�_
o
�_/o�8UFRAM%�/P!�RTOL_ABRqTSoN#kbENBto~ehGRP 1S�����Cz  A� �c�a��o�o�o�oB"v,>cj��U�h�#!�kMSK  h�ef!�kNPa%^)��%�_��e_EV�Ns`�t&�v�2�T�;
 h#!�UEVs`!td�:\event_�user\�7�C�7<�o� Fq�/�S�P5�:�spot�weldl�!CA6��r���#�t!� K�	�>��q��-�� q���Q�c�ܟ�� ��� ��ϟH��l��)�_� ����د����˯ �� D���z�%�����[��m�濑�
ϵ�Ǻ�W�RK 2U�a8�nπ� \ϥϷ� ���������#���G� Y�4�}ߏ�j߳��ߠ� �������1��B�g��y��$VARS__CONFI�V�;� FP����C�MR�b2\�;�xy� 	$ ��0�1: SC130EF2 *�	�����X�ȸp�  �#!?�p@pp:"p�z� o]�g���������������`�uA�����,� B���G�K��l�� �_������ �2�hSe��Q����IA_W�OF�]^-˶,�		�Q;%/+'G��P �> ���RT�WINURL ?5�������/��/�/�/�/�/�SI�ONTMOU� ���%�^Sۿ��S۵@�a� FR:\�#\�DATA؏  �� UD166wLOGC?  \9�EXh?'q' ?B@ ���2{1�U��?{1�?�?θ �� n6  �������2zt�`�F��  =����BA��?@|=TRACIN�?AQB�d�CpBEFF/B�0�(��_� (��I�M ��O�O�O__P_>_ t_b_|_�_�_�_�_�_.�(_GE3`�/C��
�`'p4b
g�0R�E!0a�i���LE�Xdb����1-e��/VMPHASE'  ���C ���RTD_FILT�ER 2c� �&��T��o+ =Oas�����o ������1�C��U�g��)SHIFTMENU 1d�K/
 <�<%�?ŏ2����ɏ�ُ� 8��!�n�E�W�}���������ß՟"����	LIVE/SN�A��%vsflsiv�n4���#� SETU��W�menum�r��ѯ��"��3e`+|�MO�3ftn�z��ZD��gQm˳<�A�P��$WAITDINEND8L!�k�OK  �醼 :r��S����TIM5���Gr�͔��%˴��ӿ�򿆸RELE�a5��k��/<6m�_ACTJ�4�t !��_?1 h���%�5߅���RD�IS����$X�VRnaitn�$oZABC��1jQk' ,�@�2=��-�ZIP2kQo����)���MPC?F_G 1l��l!a0L"��q�7�MP��am����P�������`�*�  4�Y��G�4/���G�Y�Ǵ��K�y5�����H�D�b���_�B��B�0�Q��5�(>����<�ȴ0+&���=I?�j�\����&?���|���&?���{� ?�.��8�}���p9��������C²��B���j�r�7�5B��³ a´ 'Gl�PJ\r� �������6��.�ȇ�J�p`n��_C_YLIND�aoR�� �p6 ,(  *o�w3l���� ��// '.iJ/�n/U/g/�/ ��/�/�///?�/�/ F?-?j?Q?�/�?�?r�Cp*� �g� �?L^���6O!OZO?Ih�?�O?G��AA�=�SPHERE 2qO�?�OT?�O_ �O:_�?�Op_�_�/�_ E_+_�_�_ o�_Y_6o Ho�_�_~o�_�o�o�o��oo�o ��ZZ�� ��