��   v��A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����UI_CO�NFIG_T � x L$NU�M_MENUS � 9* NEC�TCRECOVE�R>CCOLOR�_CRR:EXT�STAT��$T{OP>_IDXC�MEM_LIMI�R$DBGLV�L�POPUP_�MASK�zA � $DUMMwY73�ODE�
]4CFOCA ��5CPS)C��\g HAN� � �TIMEOU�P�IPESIZE �� MWIN�P�ANEMAP� s � � FAVB ?� 
$HL�7_DIQ?� q�ELEMZ�URȩ l� Ss�$7HMI�RO+\�W ADONLY�� �TOUCH�PROOMM�O#?$�ALA�R< �FILVE9W�	ENB=�%%fC 1"USE�R:)FCTN:)W�I�� I* _E�D�l"V!_TIT�L� 1"COO�RDF<#LOCK�6%�$F%�!b"EBFOR�? �"e&1
�"�%�!BA�!j ���!BG�#�!hI{NSR$IO}�7PM�X_PK�T?$IHEL�P� ME�#BLN=KC=ENAB�!? �SIPMANUA�L4"="�BEE`Y?$�=&q!EDy#�M0IP0q!�JWqD�D7�DSB�V� GTB9I�:J�<wSTYf2$Iv!q_Gv!k FKE��FHTML�_wNAM�#DIMC4|:1]ABRIGH83s oDJ7CH92%!FE�L0T_DEVICzg1&USTO_@  t @;AR$@PIDD�B�C�D*PAG� ?�hA�B�ISCREVuEF���GN��@$FLAG�@���&�1  h� 	$PWD_A�CCES� MA�8��hS:1�%)$�LABE� $	Tz jHP�3�R�}	4SUSRVI >1  < `�Rp*�R��QPRI��m� t1�PTRI�P�"m�$$CL�ASP ����a��R��R `\ S�I�	g � �iaIRT�s1	o`'2 L1���L1���R	 K,��?���aF1`�b�d~a�����y`� �`�c�o��
 �� a�o�o1CU �oz����� c�
��.�@�R�� v���������Џ�q� ��*�<�N�`�� ������̟ޟm��� &�8�J�\�n������� ��ȯگ�{��"�4� F�X�j���������Ŀ�ֿ���`TPTX��ʊ�)��� s �Ƅ��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg���Ϩ�Ⱥ��υ�&a�s�pwd���+�=�O߄�s� �ߗߩ߻���\���� �'�9�K����߁��`����������a��f�b�b�� ($p�-����T�?�x���a�a��c���c$����l��k
��a�h�ah�h�t�h�	f����������`���` � ���f qT��h#h�Fd��g��Xc�B 1)hR� \ _�� REG V�ED]���wh�olemod.h�tm�	singl�	doub �trip8browsQ�� ���u���/�/@/���dev.sl�/3� 1�,	t�/_�/;/ i/??/?�/S?e?w?8�?�?�?� H`�? �? OO$O6OHOZOlO~O�F @�?�O�O�O �O�O_�F�	�?�?;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o mooM'�o�o�o�o�o �o+=Oas �������� �?>�P�b�t������� ��Ώ���O����� L�^�_'_������� ş�����6�1�C� U�~�y�����Ư��ӯ �o���-�?�Q�c� u���������Ͽ�� ��)�;�M�_�-��� �Ͼ���������*� <�7�`�r�A�Sߨߺ� q���i�����!�J� E�W�i������� ������"��/���O� I�w������������� ��+=Oas ������� ,>Pbt���� ����//���� �^/Y/k/}/�/�/�/ �/�/�/�/?6?1?C? U?~?y?�?Y��?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __�R_d_v_�_�_ �_�_�_�_�_�o*o��_o`oro�j�$U�I_TOPMEN�U 1K`�a�R 
d��a*Q)*def�ault5_]�*level0 =* [	 �o�0��o'rtpi�o[23]�8tpst[1[x)w�9�o	�=h58�E01_l.pn�g��6menu15�y�p�13�z���z	�4���q�� ]���������̏ޏ)R r���+�=�O�a����prim=�p�age,1422,1h�����şן� ���1�C�U�g����|�class,5p�����ɯۯ�����13��*�<�N�h`�r���|�53��@����ҿ�����|�8��1�C�U�g�y�����ϯ���������"Y �`�a�o/��m!ηq�Y�w�avtyl}TfqOmf[0nl�	�Пc[164[w��5�9[x�qG���/��2 9��o�%�1���{�� m��!�����0�B� ��f�x���������O� ����,>����2P�����\ ��'9K�� ����������1��/$/6/H/Z/���|�ainedi�'ߑ/�/�/�/�/���config=s�ingle&|�wintp���/$?6? H?Z?!Z�a�h?�?�e �?�;��?�?�?OO +O=OOO�?[O�O�O�O �O�O�O�O_a�%_L_ ^_p_�_�_�_���_�_ �_ oo$o�_HoZolo ~o�o�o1o�o�o�o�o  2�oVhz� ��?���
�� .��@�d�v������� ��M�����*�<� ˏ`�r���������^��;�M�sc�_;���s��X�}���e�u��0���P��t��4�j�X�6e�u7�����ｿϿ�� �P�)�;�M�_�qσ� ϧϹ���������
�"�1�M�_�q� �ߕߠϹ�������� ��7�I�[�m��� ������������!�����6(�]�o��������$��74�������)t<ϯ\�5	�TPTX[209©|Dw24§J����w18�����02��A#��[�tv`�Rd$vL0�K1����5S:�$treev�iew3��3��&�dual=o'8?1,26,4�O/ a/s/2�/�/�/�/�/ �/�/?'?9?K?]?o?2��;/��53$/6$ ���?�?�?
?#O5OGO YOkO}OO�O�O�O�O �O�O�?�?��1�?6$�2�f_x_�_ �6<_��edit��>_ P_�_�_o��/���_ �Sooo�o�oB�o�o ��oA�o�+ =Oas��o�� �����(�9��� Q�x���������ҏ�O ����,�>�P�ߏt� ��������Ο]���� �(�:�L�^�ퟂ��� ����ʯܯk� ��$� 6�H�Z��l������� ƿؿ�y�� �2�D� V�h����Ϟϰ����� �ϕo�o��o@ߧE� c�u߇ߙ߽߬����� O����)�<�M�_�q� ���W��������� &�8���\�n������� ��E�������"4 ��Xj|���� S��0B� fx����O� �//,/>/P/�t/ �/�/�/�/�/]/�/? ?(?:?L?��߂?1� �?���?�?�?�?O $O5OGO�?SO}O�O�O �O�O�O�O�O��2_D_ V_h_z_�_�_�/�_�_ �_�_
oo�_@oRodo vo�o�o)o�o�o�o�o *�oN`r� ��7����� &��J�\�n������� ��E�ڏ����"�4� ÏX�j�|�������a? s?蟗?�sO_/�A� S�e�w���������� �����,�=�O�a� #_������ο��=� �(�:�L�^�pς�� �ϸ������� ߏ�$� 6�H�Z�l�~�ߐߴ� ����������2�D� V�h�z�������� ����
����@�R�d� v�����)����������ƚԔ*de�fault%��*level8��ٯw���? tpst[1]�	��y�tpioG[23���u����J\men�u7_l.png�_|13��5Ж{�y4�u6 ���//'/9/K/]/ ���/�/�/�/�/�/j/ �/?#?5?G?Y?k?�"�prim=|p�age,74,1�p?�?�?�?�?�?�"��6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_ �_�_�__B6o9o�Ko]ooo�o`�$U�I_USERVI�EW 1֑֑�R 
����o��o�o[m �o'9K] � ����l��� #�5��oB�T�f���� ��ŏ׏鏌���1� C�U�g�
��������� ӟ~�����v�?�Q� c�u���*�����ϯ� 󯖯�)�;�M�_�
� �~������ݿ�� �%�ȿI�[�m�ϑ� 4ϵ��������Ϩ�
� �.ߠ�i�{ߍߟ߱� T���������/��� S�e�w���Fߨ�� ��>���+�=�O��� s���������^����� '����FX�� |������ #5GY�}�� ��p���h1/ C/U/g/y//�/�/�/ �/�/�/�/?-???Q? c?/p?�?�??�?�? �?OO�?;OMO_OqO �O&O�O�O�O�O�O�? �O_ _�OD_m__�_ �_�_X_�_�_�_o!o �_EoWoio{o�o0h