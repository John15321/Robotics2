��   b�A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����CELLS�ET_T  � w$GI_S�TYSEL_P �7T  7ISO:iR4ibDiTRA��R��I_INI@; ����bU9�ARTaRSRP�NS1Q23�4567�8Q
TROB~QACKSNO ��)�7�E �S�a�o�zT2 3 4 U5 6 7 8a\wn&GINm'D�& ��)%��)4%��)0P%��)l%SN�{(�OU��!7� OPTNA�73�73.:�B<;}a6.:C<;C�K;CaI_DEC�SNA�3R�3�TRY1��4��4�PTHCN�8D�|D�INCYC@�HG�KD�TASKOK�{D�{D�7: �E�U:�Ch6�E�J�6 �C�6U�J�6O�;0U��:IATL0RHaRxbHaRBGSOLA�60�VbG�S�MAx��V��Tb@SEG�q�T��T�@REQ�d�drG�:Mf��GJO_HFAU�L�Xd�dvgAL�E� �g�c�g�cvgE�� �H�dvgNDBRx�H�dgRGAB�X�tb���CL�MLIy@  � $TYPE�SINDEXS��$$CLASS ? ���lq�����apVERS�IONix�  �i}qIRTUALi{q'61j�r���p��q̹t+ UP0 �x�Style �Select 	�  ���r�uReq. /Echo���Ack���Initiat(�p�r�
�^�m�R�����	��
��V  �������������χ�q�)��Option? bit A<��p��B��C4�Dewcis�codY���Tryout �mj�6�Path �segh�ntin5.8�Ig�ycX�:�Task OK���?�Manual _opt.r�A����B���C� d�ecsn ��$�R�obot int�erlo7�@�\� OisolQ�4�C���iM�@���ment�<�)�������Ě}�s�tatus=�	M�H Fault:<����Aler�1��C��p@r 1�z �j�;�y���I�; L�E_COMNT �?�y�    Չ�ѿ�����*� <�N�`�rυϖϨϺ� ��������&�9�J� \�n߀ߒߤ߶�����@�����"�����U���Ђ��Ŵ   ��E�NAB  �� :���������������MENU\��y��NAME ?%��(%$*R�זb�� P���t����������� ����+O:s^ p������  $6HZ�~ �������/  /Y/D/}/h/�/�/�/ �/�/�/�/?
?C?.? @?R?d?v?�?�?�?�? �?�?�?OM