��  	w^�A��*SYST�EM*��V9.1�0185 12�/11/2019� A  �����AAVM_�WRK_T  �� $EXP�OSURE  �$CAMCLB�DAT@ $PS_TRGVT��$X aH]ZgDISfWg�PgRgLENS_CENT_X��YgyORf  � $CMP_G�C_�UTNUM�APRE_MASwT_C� 	��GRV_M{$�NEW��	ST�AT_RUNAR�ES_ER�VTSCP6� aTCb32:dXSM�p&&�#END!�ORGBK!SMp��3!UPD�O�ABS; � P/ �  $P�ARA�  ����AIO_wCNV� l� �RAC�LO�M�OD_TYP@F+IR�HAL�>#�IN_OU�FA�C� gINTER�CEPfBI�I�Z@!LRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CES�0�!H1�!  � A> �1	 � �$SOFT�T�_IDBTOTA/L_EQ� Q1]@�NO`BU SPI_OINDE]uEXBSCREEN_�4�BSIG�0�O%KW@PK_FI�0	$THK�Y�GPANEhD �� DUMMY1"d�D�!U4 Q!�RG1R�
 � _$TIT1d  ��� 7Td7T� 7TP�7T55V65V75V8
5V95W05W>W�A7UPRWQ7UfW1pW1zW�1�W @V�R!SBoN_CF�!�0$!J� ; 
2�1�_CMNT�$�FLAGS]�C�HE"$Nb_O�PT�2 � ELL�SETUP � `�0HO�0 P�RZ1%{cMACR=O�bREPR�hD0�D+t@��b{�eH-M MN�B
1 �UTOB U��0 9DE7VIC4STI�0�A� P@13��`BQd�f"VAL�#ISP�_UNI�#p_D�Ov7IyFR_F �@K%D13�;A�c��C_WA?t�a�zO�FF_@N�DEL�xLF0q�A�qr�?q�p�C?��`�A�E�C#�s�AT�B�tcbMO� �sE' � [M�s���2�REV�BI�LF�!XI� %�R�  � OD�}`j�$NO`M�+��b�x�/�"u�� ����^���@Dd p �E RD_Eb���$FSSB�&W`K�BD_SE2uAG*� G�2 "_��B�� V�t:5`ׁQC�4@�a_EDu �O � C2��`�S�p�4%$l �t'$OP�@QB�qy��_OK���0, P_�C� y��dh�U �`LACI�!�a���<� FqCOMM� �0$D��ϑ�@�pX���OR BIGALwLOW� (KtD2�2�@VAR5�d!�A}#BL[@S �� ,KJqM�H`S�pZ@M_O]z����CFd XF�0GR@��M��NFLI���;@U�IRE�84�"� SgWIT=$/0_No`]S�"CF_�G�� �0WARNaMxp�d�%`LI��V`NST� CORz-rFLTR�/TRAT T�`� $ACCqS�� |X�r$ORI��.&ӧRT�`_SF\g�0CHGV0I�Ep�T��PA�I���T��1��� �� �#@a���HSDR�B��2�BJ; ��C��3�4�5*�6�7�8� �~"��x@�2 @.� TRQ��$%f��4ր����_U����zf�Oc <� �����Ȩ3�2��LL�ECM�-�MUL�TIV4�"$��A
2FS�ILDD��c� �DET_1b ; 4� STY2�b4�=@�)24����FҼ� |9$��.p��6�I`�* \��TO��E��EX�T���ї��B�ў2c2ӱE��@���1b.'�B ��G�Q� �"Q�/% �a��X�%�?sdaD�U�A Sҟ�;A�Ɨ�M�� � CՋO�! L�0a�� X�z�pAβ$JOBB���������IGO�" dӀ�����X�-' x���G�ҧ]�C�`�.�b# tӀF� �C3NG�AiBA� ϑ ��!���/1��À�0��H��R0P/p ����$
�|��BqhF]�
2J]�_RN���C`J`�e�J
?�D/5C�	�ӧ��(�@{ f�P�O3л!7% \�0RO�6�� �IT�s� NOM_8pn#�c �Ѭ�TU�@P� )� ��&+P��� bӨP�	ݭ��RAx@�n �3�A���
$TYF3%#D3
T�ԢwpU�13�}�%mH,rzT1�E� ��ޣ�#ݤ�%ߢQl�YNT�"� DBG�DE�!'D�]�P�U���@t����"��AqX��"�uTAI2s�BUFۆ;%�1( ���P&V`PI84U'mP�'M�(M�)�B �&F�'SIMQ�S�@ZKEE3PAT�zЙ8"�"԰��C��)S�0��`�JB���ľaDEC�g:� g5e�����* ��U�CHNS_E;MPͲ$G��7��_��c;�1_FYP)�TC�6S�Ѐ�5�`%��4�} ��V0����W��JR�����SEGFRAq�O��� #PT_LIN�KCPVF>���C$+���ckBZ�PB�zr�5,` + �Ԧ��A�0��Ad0�o`Ar�D���Id1SI!Zh���	T�FT�C�Z1Y�ARSm��C P@'�Ic\1@cX�0<@�L����0�VCRCߥ�sCC���U1@�X�1��2�Mpq�U�1`�X�Q�UDݤأiCk�p��
DK`݀fL��RhEVRf �Fha_	EF�0N�f�Pd1�&h��5�jC}�=+�VSCA[��AA�fK2�4��-�y	�ׇMARG��D�a�F@@���1DcQ��r�0LEW�-�@�R�P<��o�l��RɄ.� ����ǯ��� 5ڡR�`HANC��$LG5��a�� Ӑ��ـF��Ae����0RYr�3
�����
�@ �RA��
�A�Z�0Q�N`�O��F#CT��sp�F��R��0P0b ADI��O ��+���+���&���5�5����S[�g���'BMPUD(PY�1���AESCPjc��WꍠN  S-�p�C�U0ۑU�/)�T#IT'q<�b�%ECA<:!�!ERRLd�б0�&Q��OR�B$𛒿���1�$RUNs_O��SYS���4������u�REV��c�DBPXWO�P�10�$SK�o�".DBT�pT�RL�2 �C A�C����%�m�U DJ$�p�_�`�!A�ǀ�M�PL�A_2WA��j�E��D!w�!�%RhO�UMMYi9����1� �d[��3���!PR�Q�Ұ�Dٱ9��4� г$r��$ Q�Lة5�������6�z ��PC�7*�z
_�PENEC0Tq�8I�z��REC�OR$�9H �m��4$L��5$أ�"E���R@����溑_Dց� ROS �"SK�����I0�=�א��PA��J>VBETURN���S�MR(�U #�CR�ʰEWMDB0G�NALV �"$LAx� [�*6$P-��7$Pv�s�8�o�!�PC��#�D�O^@-�Ŵ���R˶G�O_AW�ܱMO�z��p��CSSW_CN4�YO�:��0T��0���ID�T�U2��2�N��O@��J��v`Iְ ;� P $>�RBl�B��PI�POl؏I_BY��vЅ�T�VR��HNDG$�< H�`�1a�@cS��DSBLI��s��h�0}�
��LS$�a=��0� ��FB��FEձL�9�����5��>D�$DO�1�C�pMC�0q��P4��9�RH��W��K4ELE�ur�����SLAVr?xBINS ���#����_R@P�@\`�p S�}�l�}�l�{u��[!"e��ے�I����B��W��D�NTV̞#�VE�$��SKAIlA4;3��2���1J�f�1C�
DSAqF7�5��_SV6��EXCLU-��NXrONL�0YY�x�s����HI_VՀ^�RPPLYo�RCs�H� �0_M�>Q�VRFY_I�.=Mms$IOv0��D}��1��Oj�F3LS����4!I��:@�P��$�ĆAUTOCNE ����.��G'CHD�s��_���36s�AF��CPe��T!��р� �Ao���_�0 s ��z�NOCtIBxB�pT��A ܢ��_SG�` �C � 
$CUR8�U��!" �� ��B�����ANNUNC�#������b���()%!��-*�I&ԢEF��IC�D� @�F
"a��POTX�aө�������l����EM��NIߢ!E�·"�G� A��$�DAY��LOAD�`Ԟ��"��5�� �EFF_AXI�%Fo�%Q�O0[��:�_RTRQV1GC D�a��?0�RK3x�0S45 2Fz@8]w:1a���A0p/1NsAH 0B!�1A�T��2�ûvDUX��u�.�CABsAIs"�p�NS�1�PID�@P�WSs�5�AWpV`�V�_�0q0�P�DIA�GysAJ� 1$VX��ET	`�UrT��EJ��{RRf��!�T�VE�� SW�|AZ�sP�0�:5q0G�}P:1OHP5�1PPL|@�SIR|�{RB�P �2�3%qZQC �BB���H�^��E`��5q0I���?0���URQDW&�EMSB�?UA�p�E<jB�TLIFE�`K#iP��uRN|QFB�U%!�zSFB�a�%"C����N��Y'p�F3LA�t& OVڰ�V�HE��BSUPPIO(��uRI�_�T��Q_X�d�� gZjWj� g��%!���6�XZ*�ϡfAY2xhC��T��DEQN�pBE%!J�� �F�_8p�A�� @C�T�K `Q�C�ACH�*r�bSI�Z�V�P`�N��U7FFI`�oP��ў�2��6���M�;��tL 81 KE�YIMAG �TM ��!�^q:�Yv�����OCVIE�@�qM �༠L~��;�C?���р�dNG0m��ST��!�r ���t���t0�t0�pEMAILo����!���5FAUL�"Op�r��/���COU���q^T��)AP<' $9�p�S�0�0;IT��BUF�g;�P�gE�o�e��PBe��p�C:���:�|�G�SAV��r�[@�b��@ˇÐ)&P��p印�D���_e���� �OT겮�3Pm ��0�zF3�AX�#f x Xe��C�_G|S
�YsN_�A��Q <�QDk�O����BM�2��PT� F�$,�DI[E7���$��R��$ G���!&�Ǳ���:�9��S����-��C	_ᰤ�K�$������RVq���DS�Pnv�PCe�IM@��\���<�3@U9�0�P�] �IP���A�`[�TH�`3�O�20T�\�HSȓ>�GBSC���`e�V���
��#���*4NV���G;���`Y�e�F�|A}�d>���Z��SqC%Ba��MER)>�FBCMP)��ET�� TLrFU`DUY���R�mb�CDR�ܠ'�"���QR��n!UG0*А���%���%P���C"�
ō-"2��|:�o VH *
�L��)�9���G �� ��}�Z{ƥ!{�1{�P1{�6q{�7x�8xɡ9x�|PzȄ�1��1���1��1��1��1���1��1��2��2T�ˑ�2��2��2��U2��2��2��2�ʕ3��3��3�˞�3���3��3��3��3���3��4��61EX	T6An!W��߸���V���uş�����F{DR%DXTE��V� .�uR�
�uRR�EM^@F���BOV�M5�*�A3�TRO�V3�DT��S�MX�b�IN3��PR�"AINDq�cB
��ɐ}���Ge��C\�p�UkA9DO6\�RIVW�R��BGEAR5�IObEK#�cDN��1�`X� zp`dCZ_MsCMp`uQ��F�P;UR��Y ,����? �P>?\o {A?oE� w��*�������Z0*PPM�2@R�I��0r�ETUP?2_ [ 0q�#TDʠ�1p�T��p���1r�BAC��G\ T�pr��)��%w#@ó�TIFI��A����d��@/PT��B�qFLUI�t�] �@�x;�UR �A���R�Б
��:C�_0I�$�S_k?x�J�CO���"�VRT��� x$�SHO^14 #�AS�S�-��U̠��BG_ �!.�!��!��<!��FORC�i�DATA)A^�rF%UZ1��]#2��5��i�`)A_ |��N;AV=�������S��S$VgISI��SC=��SE� ��5V� O
�1&1BF�4@�&�$PO� I�A��FMR2��` ���2� ��6�!3J�)��CE#�_����_@I#T_Yִ]@M�������DGCLF�ED7GDY�8LD���5�V���T��0�ua�4�v9 T�F9S
��tb P��RB|��}�$EX_RA�iHRA1Y�X��RS@3��K5�F�G&�	5c� ���SW��O>0VDEBUG$�A�(�GR� opUz�B�KU��O1M� �0POZ0Y�@��t�E�@M�LOOM�9QSM�0E��J�����P_E d �rp��TERM[Ue�dV�pORI֑`PfdU��SM_��`P�g}YQ �XhdU��U}P�ri� -��F�2d�rS�Pe� yG�Z @ELTO�9��A�FIG�b�Z �Agp�T�Tf$U;FR�$��a�M`ѵ�0OTZgA�TqA��lcNSTא�PAT��`�bPTHJ�ϰE�p�ذbART؀"e)�؁����REL�j�S�HFTӢ�a�h_��R��̳�V �P$�Wph�1����t��SHI�`�4U � ҁAYLO��m����l� ��a}!�ޠERV��Sq�x��hg�א�b �K�u.�KRyC��ASYM����WJ+g���E ��a�y�ұU�א ���e@�v�eP��pp�E�2vORאM3��@JQ
4jX"�B0V0�`G`l�� HO�6D�k ��aN� �O�CaQ@$�OP�$e�i��H����ՀRY���aOU��c�PT�R�e����ae$7PWR��IM��rR_˃�d� �P�c�UD��cSV��t��֔l� $H畽!��ADDR��H�MQG�b������L�R\�"1m H��S�� �! ��.�畞�畫�cSEz1�#��HSܰ�
3n $� À_�D��P�.�PRM�_�"t!HTTPu_��H1o (���OBJ� ��$���LEyc��d�p� � �睱AB%_��T@S��S����{KRLK�HITCOU� À�!퀀������M�S�S��v�JQUER�Y_FLA!a��B_WEBSOC�"G�HW��a1q�}7�INCPU�B�!Ou�ˡ�Č�����������T�IOL]Nr 8��R	ި $SL2$�INPUT_PQ�$�ܸP�#r ��S�LA�1 sð�ٿ���s��r�QI�OC�F_AS8Bt$L&��&q�!]�/a�ɳ�@ҳUpHY���l�UQG�wUOP5Eu `X� �����ā������P�����������pC¬�qqv l�@�;sTAkr��A�T�I��.�a�Z0S��`PmSR�BUZ0ID~0 ��z���yը  �u�&z`w�3�f�G���N��Z0���IR�CA��� x �Ĩ��CY�EA{���!���%�¦R�`�q|�8�DA�Y_��}�NTVA����i�¦eu�i�S3CAepi�CL���"����� qy����X�b����N_ՀCQ�Ђ�W�rz�O � �������y�G�]�O!? 2y ��"фq{P���P�L�ABzan�Z0t�UN�ISb�PITY0��"ѳ��QIR$6D�|R_URLޏ �$AL10EN��@�� �PH�T�T;_U� �Jt�q} X��t�R��" �0A�D�,J�8FLt@�80�
K�3
�UJR.	5~ ���F|@1w��FgwD��$J�72�O!�$J8B�	7�@\��7s�� 8�	�APHI�@Q��Df@J�7J8�
L_K�E��  �K���LM��  �<��XRK��� �WATCH_VA�!�pp��FIELDb��yu &��� �0bpaVyp�ֆCT����E��B
��LG~���� !��?LG_SIZ���@`�3@�O��FD�I��,Q��]P� ���J&3@J&O�J& �J&]PJ&�q�E`1_CM^c�!{@�*h1AF��'�$��(�#r��&3@�&O��&��'I�(�(,P0�&]P�&�RSI�`o  (�PLN�
�B�����@{A�@g1��K�u1��L~3nt2DAU�5EAS�0�����2�0GH���Q�[�BOOܑ�g� Cr�[�IT8���4<`n�RE(��8ScCR� ڣs�DImùSG`G@RGIPR$D/L�f�քYB��[�	S��Z�W7D[��4f��JGM�GMNCHLH�[�FN�FK�G���IUF�H2p�HF�WD�HHL�ISTP�JV�H�P�H�0�H�RS3YHJ��Kc�C�4tS�f�x�kG�YU J��DjG 3yE�{��BG�I�`PO�WZ&E�S�"�DOC���FE]Xb�TUI�EI/  ���/!�dDa�CNc�@��p�� 4	��EpvANOGfANA[�ā�AIt瑜��DCSZ���c���bO�hO�gS?��b�h9S�hNHIGN���`��A�(��dDE��pTLL�q��|A��*�i����T�"$����}��Ԫ�SA������ʰ��Z�� *�P1�u2�u3�q`�8br�a*І ���V��c��5�z�x�6���P�6�.�ST��R�0Yy��`Q� �$E_�C_�� I��n�����T)ч L o���瀖�x������_�ENS�_�ppBC/_ �����X�x��@��MCh2�� ���CLD�P��TRQLIp��D�2�FLGZ�2�3�f���Duf�`��LDf�P�f�ORG�jQy��(RESE�RV��Ŕ��Ŕ��#�3�� � 	0O�jUA�f�SVX0D��R	���'�RCLMC5�şןG���D'�M�MՠJ�/�3�$DEBUGM�AS��S�D�"��T԰`p�E� TZ�
��MFRQ��� �� �HRS_KRU�ځ�A)���UFREQ� 8�y$``�OVERh�����v|P�AEFI��%�������9�ѣ� \ �ν$U��?�����PS�p7 	��C�06�BҒ�G�U|�Н�?( 	��MISCi� d�q1�RQ5		TBB@�� ��aa��AX9�!	�"�EXGCES��"ܲM��
.����9�oܲ�SC� � H���_G���,��� �2�ڰK���|��B@���B_�FLIC���B@QUIRExSMO��O��d��0�ML܀M��� @
��19Э��5�`pGMND�1e�/�o2�f2�x�D�#�4IN�AUT(A�4RSM� ��pNZ�b!�S^�{�d�PSTL.w� 4��LOC��RI1P�EX��A�NG�b��ٱODAե��p�x MF�%7�+�ۂ|@p�e�c0��SUP�v�pFX/ IGG�1 � ���ۃb! Cۃ�Vۄ��V�P��� R���R�����SD�w���TIj�p�pI�N��� t-�MD*��)8��`C�L�@�qH�C�DIA�D�2 W]AC��q��C�-D�3)�m�Oh�n/� a�CU��V����q�OPA_��.� �/��7�L��f��
 ��P��h>P���P��KE�RR�#-$B������ND2N�ND2_{TX�XTRA�c4p`��9�LO�0/��_���i2�����1MRR2>൜� -��1�A$� d$CA�LI��c%G�a�2ξpRIN�!�<$R� SW0S� `�wABC>�D_JV �����7�_J3K
�E1SP���P�El3k�񱀦�B�J`����Oiq�IM`�ŲCSKP S��� �c�J�1Ų�Q�%�%'�_cAZ#��=!ELNq<�N�OCMP�Ʊ���z0RT��h#�11����1��(o`:�*Z�$SMGMP�vn�JG�SCLB���SPH_�`Ű+0��#\ ��� RTEIR��`� _�`
�*�AP@G�Ų4sDIS!�"23U�kDF��<1LWB87VELD�IN�Z`e0_BL�`��m4����J]4r7�7�4��IN� ������5QBҦ���1��_̰ ���5�2#5�3�1z�936N�DHB�r ����p$V� ���#�oa$� �����$\q�R������H �$BEL�N ��!_ACCE�s1 �H`��@IR�C_0���NT<��/�$PSB�7�L����DL��0�G 3�`�F;�I�G�C�G3�B��E�_�qPB-Pp3Q����A_MG��cDDPQ2��FW�����ClU�C�BaXDE��[PPABN�GRO� EECR�q�_D��!�q�����A��$OUSE_� �cP�CTR�dY�Pb@"�- ��YN߰Aa`f�Z�aM����bJPqO_0�AGdINC���RpT�ig��ENC0L��A�B,��@IN7�I�B�e���$NT]3�5NT�23_@2���cLOQ0���`-�IP����f�F0����� ���e��C<�0�fMOSIUQ�����3Q�ŲPERCGH  s+�2 ]w �hs��rn���c'["�e
P2P�A�B�uL �T�����e��z�v�vTRK�%ʁAY ��s��,��B;�0��pn&��wbȠMOM��»������S�0G��C�R� DU�(R�S_BCKLSH_C�r����<v,�"c���݃�b�1a%CLALM�d��m�@��CHK��NGLRTY��5�d���r�_Z�1t_UM���l�C��^Q�!����LMTh_L��V#��j�E��Ð�����E����H}���r��xP	Cnq�xH���TUl��CMCv^PbWCN�_�Nuc��SFtA�yVb�g�!8���r��<�CATs�SHZ��bT�f]����f`��A�	� QPPAs�&gb_Pr�V�_�� �3�Qp�C�U�F�JG0>�X�I�K0OGV�2TORQU�P�/s�L��P��Gr1�P��_W��,��!QAٴBCصTHCصI�I�IHC�F$�˱�-��ZPVEC�@0����N�1T�pRPh�$!Z�JRKT�X�ƴ�DB� M��:��M��_DLBA�rGRVߴ��BC��HC���H_����@�CcOS�p �LN�� 6�W�=�B@8ٵ 8�
�t�b�(���Z1�Gv��MY?Ѳ��='����THET0uNK�23HC��<C@�CB��CB<CC� AS��'�
�5�BC5��SqBBCS��GTS��QCo/��'��'��q�$DUC��w��P�t5��5Q�q_�V�NE��AKS�z)!8 @��A���'�8���LPH����e��SW�o�b�o�q�@��֙�����V@�QV5�2@X�Vg�Vt�UV��V��V��V��V��H@�Y�_W�ܡTvt�H��H��H��UH��H��O1�O@��O�	V�Og�Ot�O���O��O��O��O��F��"�~bՃ3��SPBALANC�E_�ѮLEj�H_��SP�1S��b�|�q�PFULC�`"�"q��:1�|!�UTO_>�F�T13T2B)�B2N%��B �`b$�!f� ���B}C���T�pO50�AɰI�NSEG�B qREqV�& p�aDIF�f�91��'321��COB�!	��Ó�2����`0���LCHWA�R�R7BAB%���$MECH+���9a,?1T�AX9�P�X68�#B7 � 
Y2���{A�eROBQpCR��r�5M�T�C�yA_A�T � �x $WEIGH6`�$1��3X��I6a�`IF�QjPLAG'b�S'b� 'b7BILEODo�#p&�2ST�@�2P�!	�B�0 `@Ơ�1�0��0�
�`yB(aA�  2y�.t�6DEBU�3�L�@<B��MMY�9�E� N��D�3$D�Axq$�@S���� �D�O_�@A�1� <@�0VFL U�(a�B&B@N�c�H_p(`BC�O� �� E%��T�`�a��T�!<~D�@TICK�30�T1�@%NS��WPNQp1 �CQpRԀ(a!2�iU!2uU�@PROM�P6cE� $IR��&aL��R�p�R�MAI��aa8b�U_�@�S� B�:`Rn��COD[CFU.`�6ID_ppe� �R~�G_SUFF
�G Ca�QdR�DOlW� mU @lVGRC!2Id�SUd!2`e@!2le��Id�De@��0�H� _FIZA9n�cORD&A �0��B36��b&a�@o$ZDTe	 BB��E�4 *�!L�_NAQWPriUDEF_I)xr�V5t uU-BhV7DhVasuUou�VIS�����A��hTD�suS3t���D4l����7BD5 ���t[CD�O��BLOCKE�Cci_{_�W�qIbC`UMHerIdasId ouId�rUbK�TeDsUd tUb5F���q`c,0B� `er`eas`c���EhPP� �t,P�q��@�W*�)� � ��TE��D�� ALOMB_tC�^�0�2VIS!�WITY�2AS�O'CA_FRI2#��� #SI�q���RTP���_P��3tC�2W��W���������_��jaEAS�3jbd������pT�R��4��5��6�3�ORMULA_I���G	w� h� �N7�ECOEFF_O;Q� ��;Q�r�G��3S�0�BCaA �O�CCAGR��� � � $h �u"�BX+PTM��� �AR(�%��CER�� T	�te@�  �+"LLkd�pS�_3SV�tw�$L�e@q���v�e@� ���SETU�sMEA��P(`F��0CA�b�0�� � ���0  �@o��Q2��q�r�WP�q��tբ ܑubÕQ�p�q�p�+���� �PRECt�a�qSK_���� P�11_USER^!N�}�08��}�^!VEL"�}��0��!1I�`J ��MTQCFGs��O  YP� OG2�NORE�0P����0��� 4 pݳB7�2H1XYZ�c�J!o yCH0���_ERR�1� �I�Q��Pۣ@�aAi�����@BUFINDX����o MOR� H�0CU@�QH1����Q�a���"�a${0��~q£0�;���G� � $SIj����P�!Ɓ�VO����0OB�JE���ADJU�B�� �AY�p5��D.�OU�`Վ�'a.�b=��T� ]�8��\��BDIRa�i�p� ��"�0DYN�$�2��T6 �R��,P�&@��OPWOR��� �,�@S�YSBU �SO!P��cҎ���U��� 1P ����PA���X�C2�OP^`U�!���!XB�AI�IM�AGS��0U�7BIM��o�IN��@�n�?RGOVRD��	���K�PM�m�0� ߀(�s��H2L�B=з >�PMC_E�`cъ�ANM��A�B1��BP��SL�t��{ ��0OVSL�&S�DEX�q}p/2G2� ��_��G�` ��G�`Qfa�B��C�0p�%�c��_ZER����s�G� @вb5O`RI��s0
��P�	���*l�PL��Ĵ  $FWREE��E��H�T� �Ls����TD0�;@ATUS㰤AC#_T��r�UB�_�H��s�A4�`t��C D�AI�2RL���a2S�an S���XE@Y������ ��0XUP��p�qP!X�PF�D3�����PG�Ÿ��$SUBGb5��G��JMPWAIT8�V_%LOW�BQ��@CVF�QZPG2bb!Rz���U3CC� �R��MR�'IGNR�_PL�DBTB2;@P�qH1BW�P�$2��UP�%IG0�P=IG3TNLN�&2�R�����N�P)P�EED�8HADCOW;@�����E7pS4F1!4pSPDs�� L�0AV�5ps0�3UN�0"+0!R��LY�`� QN���P��v1�G�C$��M�P�@L+.�NPA�T�2xDN��PIP%w0���ARSIZ�T��c�|q�Om`�h�AT�T���"\�B$�MEaM�B�A>C�3UX��̬��PL`�ļ �$���SWITCiHZ"�AW��AS��i2�BLLBv1�� $BAZ�9D�s�BAM� ��4�I��@J50�����B6�F�A_KNO�W�3R��U!�AD��H۠~0D��5YPA�YLOA鱱�SS_Ps�\W��\WZYSL��yA�mpLCL_�� !���R�A��T�T���VF�YCK�P�Z貓T��I�XRM�H�W_ҬTB���J)�a_J�Q����AND^�9�8d�R�Q8���PL�@AL_ ��@~0���A��k��C"�DXSE!��J�3M`af� T��P�DCK��r�CO>Ű_ALPHqc�c�BE��W�qo�l	��Т�!�� � �\40R_D_1YZ2�TDŰAR�4x!uEv�0s��TIA4_y5:_y6"�MOM��ks��sxs�s�s��Bv A�Dks�vxs�v�sPUB��R�t�uxs�u�r�}Fp��� L$PI�1s��^W.���xY.�I:�IH�I V�<p}Q7��!�� !���b�ӆ��73HIG�C73w%p4Іp4 w%� z�І�߈�!�<�!w%SAMP����B�ЇC�w%�@>c 5�q���7 �Ҁ�  ��p0"p��0p������`hp���	���INќ �&�ؘ��ϔw"ښ�x��:�GAMMƕ�S[%�$GETH��o��D�d��
ϡ�IB��2I0�$H�I�_��sЩү�Eĵм�A��٠ʦLW �����٩�ʦ�b��t0caC�%CHK��4� 	��nI_%��� ��\bxΑ�����s����v���c �$^�h 1���I� RCH_D��'� �$)�LE��������hذ�0MSWFuL�$M�`SCR
(#75_����3��d� ����kp��x�p0��D;SVv1�P��v��Kǿ�	���S_SA��A�����NO�`C ���d����d_v_ \�J�:ۂ�+R��w�0sD<�4���40��zʴ� ʈ��چ�1����Օ�ԙS�A�M�� 7� ��YL,�a������-���-�� ��b��9�az�K����W�{����py�Ȳ�M� ��P��`a��$ 7��"�M���� � $����$W���ANG ]�Q���d���d���d��d� נNP���C���ϐX�0O�cΑZpq��� �� �<�OM��"��1�C�8U�g�bpCON��0�|���a_�B� | �a�����y7xs7�s ��dzdO~z�A���4�����0�PP� A�PMON_Q}UG� � 8�0�QCOU��ǀQT�H� HO&�� HY�SD@ES�B� UE�� ��@O5$�  �@P�৥��RUN�ZY�0 O��� � POP+�%���2ROGRA��x@:�e2�Ov+IT��xINFO���C �A_�8���1�OI�� (ʰSLEQ������b=_S_EDd � '� ���r�K�QI#5��EȠNU'(�AUT��%COPAY�Q��8,���M���NB F+U�PRUTZ� I"NF2U�B�$G0�$�aPR�GADJ!�BX_��2$�0�&~�
�&W�(P�(��&73�� �NH`_CYCz���RGNSDs���LGOb���`NYQ_FREQ�rW����^1RD)L�P:BV0�!�s����CRE���c�IFlH�jNAK�%�4�_G�STATUx å�MAILI��S&@V��ǀLAS�T�1�a04ELEM�:1� �EaNAB<�0EASI&A�� v�n�?�B���GF�����I���U2����� �|BAB�C	PRS�LV	A�Fa�I��b�qU����JP'c~�FRMS_TRvC Α��Ci����A�DXXa13��& 	SB? 2�  �V� �9V(b8WR��RNTdW&�
�DO�P�W}�L�04PR �;0���GRID}�BARS��TY'C�ἐ�O�p!� _"�4!� �R�TOo�74�� � |� P�ORXc�	bSReV�0)(d fDI��T!pAaTd��^g��^gQ4\i[�^g6\i7\iI8@a�Fj�:1�?$VALU�C���9D� F65��C !"E��l�S�1���_@AN���b�1R� c17ATOTALXH��qCsPWK3I�Q>YtREGENWzlr�X�H@c5v� cTR�C�Wq_S���wlp\CV�!���u���1GRE5C�P�6B�+.  sV_H�PDqA���p�S_YѴi�o6SV�AR��2�� �"IG_S!E�3�p b�5_/�t{C_�V$CMP����DE�M���IBe�Z��^����F��HANC�� �p&Q$E�2���I#NT?`iq��F%��MASK=��@OVR�P� �P��1Α�W!a�T� 4�� �_XF�{�V�PSsLGV�:1� @K@��p5a���ApJpSh��4��U>�!��sTEa��`���`��U�Jd���3IL�_M~4���p� T�Q� ����@-�\�V�4�CB�P{�4AL�M�c�V1b�V1p�2��2p�3�3p�4�4p����p:����p���j�|�IN�VIAB��<�)���0�2,�U28�3,�38�4,�!48� hR�S��� ��T $MC�_F�  ���LP����ׅ7pM8�I׃���S ( ��n��KEEP_HNA�DD��!ﴙ@��C��0��Q��?��O��| ���p�܇.�REM'��IqPbL�c�h�U�4e��HPWD  ��SBM��PCOLLAB��p��5q�2�IT50`�w"{NO��FCAL�ܔ��� ,��FL|�A$SYN����M� Cq��XpU_P_DLY!��DELA?�Jq�2Y֨ AD��QQSwKIP�� �`-O;�NT�]�i�P_-V��^U�*� ���q���q��u`�ڂ` �ڏ`�ڜ`�ک`�ڶ`z��9wA�J2R0Z� �L�EX�@TX3 N�7AN� �N�}��`RDC��� u���Rz�TOR� ���R�1�����;TRGEA�rh@��R�FLG�^�5�ER����SPC�1U�M_N��2TH2�N�Q�A� 1�  �A��Q62 � DKш�鞝@2_PC3]�S����1_0L10_C�}2�1��� �� $b� ��� 	ViR����0�� �\Ub����mrj���C�a2��=��IDr� Gy�XUVL1a��1n��� 10c�_�DS�������P�11!� l�����#C��ATE��$�Q ���f��;T��3�HOME� )�h2n�t�������3n��'9K�4n�n�����W 2f5n��`�/!/3/E/ e6n�h/z/�/�/�/�/�7n��/�/	?�?-???c�f8n��b?t?�?�?�?�? �fS���!�.�p�Ag�p��
$C1�ze�Ed� TC�tD:vtCIOꑔIIt@f�O��_OP�EиC4r��;�R� WE�� ^@�l�8d�1�4t ���B�$DSB��GNA���3s:�C��`�QR�S232zE� ����5���ICE;US=sSPE(��a�PARIT �2qO�PB���bFLOWFO�TR9@?rt�UX��CUuP���aUXT���a�ERFACtZTT�U.p���wSCHa� t�b��_`Py���$ �&�pOM8���A�������UPDư��q3PTU@��EX��#hc�EFA8������RSP�P�a��|�`�7$USA�X��9��EX�PI��$(`�pY�eR_$�q�`mQ�fWR�OI�D���f��FFRI�END��L�$U�FRAMc�pTO;OLvMYH��r�LENGTH_V�TE�dI�;s��$Z pJxUFIN�V_^ ��_ARGuI%���ITI��bBwX�Sw�vG2�gG1�aꀎc�r�w�_r�O_XP��L�+q4���N�Sc��Cp�Pr�q�	�G���Rǁ󐒧�XQ؂��h�U���U��,�����PUd�X nm`E_MG`CT�c�H��h���U�dScG��W�`ć��لD]и@KȅJӂй�������$-� 2!���an �i1�h�`U2�k2=�3�k3�j -����iK���F�`l�P�`x�|�NtV�uV�ТPq,��r�P��� �V������R��pr�.���E9�<�Os�)E$A��T�P!Rh�U�k�ǓS��P����Sb;Q� ! �ႃ"��K��"����S`�p�p��
��$$C��S��[���P��9�9�� ؠVERSIܧ`���i��I#PP��AoAVM_�a2 �� ?0  �5�V�rb�S��� ��A	a ����9� �����ζ����ϧ�`�R�d�l�0�BS^ �r1�� <@ϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G Yk}����|»CC`XLM�@v����  d��IN����qEX$?��2_`=�r ���0�IOCip,q ��PZXQ���{�IO'PV �1=�P $-��`ұ�!̺ �?�� � ��//%/7/I/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�O__ +_=_O_a_s_�_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�o�o�o�o �o�o�o#5GY k}������ ���1�C�U�g�y� ��������ӏ���	� �-�?�Q�c�u����� ����ϟ����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i��{ύϟϱ���� LA�RMRECOV �I��LM_DG �����_IF ���p߂ߔߦ߀��^���������, 
 �G���@�m�����$_� ������ �2�D�V��h��NGTOL � I 	 A�   ����� PPINFO %� $������  1�I
�8 r\������� &W�p�Rd v��������//*/x�PPLI�CATION ?}����LR Ha�ndlingTo�ol y" 
V�9.10P/25���5'
8834�0z#�*F0�!�/1�31y#�,�/�"7�DF1� 5,y#No�ne5+FRA�5/ 6�-B&_�ACTIVE�� � [#��  X3U_TOMODb0)����U5CHGAPO�NL�? �3OUPLED 1M�� �0�?�?�?O;�CUREQ 1	�M�  TIL�L	XOiE_ ~D�wB�m%�MDH6E�2cJH�TTHKYwO��D\COUO_�O7O�O __'_9_K_]_o_�_ �_�_�_�_�_�_oo #o5oGoYoko}o�o�o �o�o�o�o1 CUgy���� ���	��-�?�Q� c�u�����󏽏Ϗ� ����)�;�M�_�q� �����˟ݟ��� �%�7�I�[�m���� 믵�ǯٯ�����!� 3�E�W�i�{���翱� ÿտ�����/�A� S�e�wω��ϭϿ��� ������+�=�O�a� s߅��ߩ߻������߀��'�9�K�CET�O��d?X2DO_CLEAN�?V4���NM  �� O*�<�N�`�r�NDSPDRYR��&U5HI�0�@��� ��&8J\n�����R8MAX@I ��|�~A�7�X����!�2�!X2PLUG�G�0���3t5PRC*��B������.O3����SEGF�0Kz�������//&/^�LAP����Cz/�/�/ �/�/�/�/�/
??.?�@?R?�3TOTAL���3USENU
��; ��?~B@�RGDISPMM�C��AC��@I@���4O������3_STRING� 1
�;
�kM�0ST:
)A�_ITEM13F  nT=OOaOsO�O�O �O�O�O�O�O__'_�9_K_]_o_�_�_�_�I/O SIG�NAL-ETr�yout Mod�e4EInp�PS�imulated�8AOut�\�OVERR�� =� 1007BIn� cycl�U8A�Prog Abo�rc8A�TSta�tus6C	Hea�rtbeat2GMH Faulug~cAler�i�_�o �o�o�o�o $6H ��/K��AO K������� �)�;�M�_�q�����৏��ˏݏ_WOR �/K���=�O�a� s���������͟ߟ� ��'�9�K�]�o�����PO-Kia��-� ��ܯ� ��$�6�H� Z�l�~�������ƿؿ����� �2ϴ�DEV��]�ЯJτϖϨ� ����������&�8� J�\�n߀ߒߤ߶���>��PALTu}� -���)�;�M�_�q�� �������������%�7�I�[�m���GRI� /K�������� ��'9K]o �����������0Ru}I��# q������� //%/7/I/[/m//�/�/�/7PREG �� a�/?'?9?K? ]?o?�?�?�?�?�?�? �?�?O#O5OGOYO�]��$ARG_�D ?	����A��  �	$�V	[��H]�G��W�I�@S�BN_CONFIQG�P�K�Q�RQ��ACII_SAVE  �TQS�@�TCELLSET�UP �J%  OME_IO�]��\%MOV_H8VPi_o_REPL�_��JUTOBACK�AQ�IQF�RA:\�+ X�_�&P'`T`�'�h� k
P �18/02�/09 11:0/6:04�&�H�-`{o�o�o�o�\���o�%7I[�&� �o������n ��+�=�O�a�s�� ������͏ߏ�|���'�9�K�]�o���X��  �Q_�S_\A�TBCKCTL.TM����ҟ����.�[INI�AeV~�SMESSAG!P�/�Q�@SQD�ODGE_D[P$VUb��O_�q��SPAUS�͠ !��K ,,		��@�Eѯ ߧů������Y� C�}�g�y�����׿���ӿ�������TSK  ��o��P�UPDTh�-�d�~�~�XWZD_E�NB-��J��STAp,��A~ŎAXIS�@?UNT 2�EQ�P� 	D�
�V���5�� �$zӟ9 ֘Y�*�� E �ASXjE�!*��=�O������@~� ��$ �~9Bv 2�r,�RU�%2hp6߿߉F��METK�24�-S P��B��>B���C�
AH>l�ZB�M�B�K���@@4?6���?�]>]0��?Lc@@�����SCRDCFG� 1�E�Q �)UR�߆��@�������o�*Q%Y s�0�B�T�f�x����� ���������,0�����G�QGR��r�X��k��NA�P�Ks	�Th_ED+��1V�� 
 ��%-��EDT- Y�Z�M�
TzPQ-�S��*�B�oxtV��  ��u2~�[\���'�@/Yk/�w3J/ ��/��s/�/%/7/�/[/w4?�/c?�/ �??�?�/?�?'?w5�?R?/Ov?�OvO �?�?eO�?w6�OO �OBO��OB_�O�O1_�Ow7z_�O�__���_oU_g_�_�_w8Fo��o��oo�o !o3o�oWow9�o_�o��;��o�o�#wCR}�_*� <��]�p���_���k � NO_DEL�w�GE_UNU�SEu�IGAL�LOW 1�	�   (*S�YSTEM+�	�$SERV_GR���*���REG3�q$U�Q�*�NUMX�<}�k�PMUրQ՟LAY��Q�PMPAL,�>��CYC10��ʞ������ULSU`��l�̒��5�L�~?�BOXORI\��CUR_,�k�PoMCNV��,��10����T4DL�I��%�G�	*PR�OGRA2�P�G_MI�����AQL¥����B��*�$FLUI_RESUЗX�b�����������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��1�C�U�g�yߋ߀�߯�������H�k L�AL_OUT ��T�WD_A�BORѐ��jO�I�TR_RTN  �st��O�NONgSTO� z� b��CE_RIA_IL��z������FCFG �
t��s}��_PA9��GP 1����Q>�P�b�!�IC�p����z�C��C ��(����C8ʅ�@��H�� CX���`��h��p��x�}�����𰂅�����	su?퀫�HE��ONFqI��Y�3G_Pr�1�� ��ă� }��������3KPAUSI�1`�� ���C `1oU��� ����/5//Y/�k/Q/�/Mo�NF�O 1`>�� � 	-��/��p� ��B�vſ��X��n²�C~�������	����	(>B��hC�3��9!C�2��1��@��D"(>�N���a�3�]گ�2����O�����sw�COLL�ECT_���&A���~7EN z��ܚ2W1NDE�3�7eヂ1234567890�7�~rD����?�6ss
 ���q)9O^OD�8O JO�OE�|O�O�O�O�O �O/_�O__w_B_T_ f_�_�_�_�_o�_�_ �_Ooo,o>o�oboto`�o�o�o�6B�2�;� �=�2IO  �9�1yxy�as؅�/wTR�2!}�� Jy
�o�~> �">}�z���9_MkORr#
� �'	 X��!X�p�^�������P��1� �q$?�,CI?,,��UpK�(TqJr��P[2&�?"�A+�a�s�����
R���t7���u�y���85���s ���9�PDB/�(7��dcpmidbg��]�v o�:��nD�p�I���m�  �b�nG�毱��ï؏�.�����mg�x�C�Ůfg����-|ſ�`ud1:����z'�DEF Y'y(Is)��c�buf.txtϸg��%�_MC8�)D7�!sd�ō�7�*���������|�Cz  �B3A� D��C����C-y�CWZ�Џ����-�Ed�1E����E9KD����E;�#��-G����G�?kGW�6�F�NGW?eG��|ɰ�(Vq���,|��t7�AUpH b�H ޒH ��t
��� ќ�@ Da  D��  E	� D��@ ���-F| �Fp F"� �G=�fF���G'i;�>��Gg� GK  �H�<=H�&�HyMc��  �>�33  `C�/��n)���5Y�T娂��A�|�=L��<#� �Vq�����ξ��RSMOFST %8ʝ/�&�P_T1��DE ;-3����q��Tq;������??���<�;��EST2�+8�PRb�2.a?����C4��%�|��Up���������C��B���C�����H�Up:d�� ���T_2�PROOG ���%x��V$INUSER�  �5($KEY_TBL  ��"�	
��� !"#$%&�'()*+,-.�/�7:;<=>?�@ABC2�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������0��͓���������������������������������耇�������������������s��q* LCKtx��&t STAT����_AUTO_D�O�6���IND��4�}1R���T927/�STO@/� TRL, LET�E�7~*_SCR�EEN ?�_kcsc�2Uo �MMENU 1/.� <ED? [�/?J?ճ'?M?�? ]?o?�?�?�?�?�?�? O:OO#OpOGOYO�O }O�O�O�O�O�O$_�O _Z_1_C_i_�_y_�_ �_�_�_o�_�_oVo -o?o�ocouo�o�o�o �o
�o�o@)v M_������ �*���9�r�I�[� �����ޏ��Ǐ�&� ���\�3�E���i�{����ڟ��ß�Ϲ�#_?MANUALs/�!�DBCO RIG��'�/�_ERRL&2 0��a�N���쵯ǯ P�NUM�LI;�Z!v�d��
�P�PXWORK 11����'�9�K��]�o��DBTB_��! 2��ç�����DB_AW�AYX�a�GCP� ��=E�ö_AL;��òT�Yr �%��I�_r� 13#� , 
�T��B�,ω�_M I��Ѽ�@����ONTIM6�'��������
�$�MOTNE�N��z$�RECO�RD 19�� y��ψ�G�O�O� =߈�Ҳ{ߍߟ߱�H� ����O��s�(�:�L� ���߂��ߦ������ �� ���$���H���l� ~��������5���Y�  2D��h��� ������U
y �Rdv��� �?�//*/� N/9/G/�/��/�/�/ ;/�/�/q/&?�/J?\? n??}?�??�?7?����OO�?9O$O �?oO�?�O�O�O&O�O �O\O_�O5_G_Y_�O�ZòTOLERE�NCдB��ްL���P�CSS_C�NSTCY 2:J����i_���_ �_�_oo'o9oKoao oo�o�o�o�o�o�o�o��o#�TDEVI�CE 2;�[ ��vu���������*��ϭSHNDGD <�[��Cz|{�TLS 2=]}<�����Џ�����>��RPA?RAM >0� ���|��}�SLAVE� ?]�I�_CF�G @J�*�d�MC:\�PL%04d.CSV)�b�cџ�RA ��CH�o�o�*��F��w�76��1s�a�<�1�JP��3|�頪�r�_CRC_OUT A]}���.�_NOCOD�~�B0���SGN� C&��&j���21-AP�R-21 01:�24�*�09�-FEB-18 �11:06��v? LIX�v�r��*�s�Iu5�M���Þ���������VERS�ION -��V4.2.10���EFLOGIC� 1D�[ 	��8+�ɘ�!��PROG_ENB�\e�A�ULS�� d���_ACCLI�M���������WRSTJNT0���*��MOJ������INIT �E�Z&�*� ��O;PTy� ?	�����
 	R57Y5*�+�740�61إ71�5�[�1U�2�1��8���TO C ݉����V���DEX��d��Hp~��PATH ۦ��A\��9�K�[�HCP_CLNT�ID ?Ѷ�� ��? ��RIA�G_GRP 2Jޣ� Q �	 @K�@�G�?���?l��>���@�����Q ����ᴝP|)��?�b�?P�T�i�^?�Vm�?Sݘ��f�403 6789?012345{������� ��s���@nȴ@i�#�@d�/@_�w�@Z~�@U/�@O�@I��@D(����@Š��p����PA�P�P�B4��Pjp��ط�
��1���-@)hs@�$��@ bN@���@�����@�D@+����������	 ���R��@N�@I�@D��@>�y@9���@4� .v�@(?��@"�\Pb�t��L�@�Gl�@BJ@�<z�@6��0��`@*� $N��@��� �$=q@����F@|��@33@�R�@-?����?��`?�+ hz����Y"J��-@&�@�N���!?�?� �� //*/</�-�/? �/&?8?�/?Z?�?^? �?�?@?R?�?�?O�? 4OFO�?VO����9 �Q�i @��V�A�Y����?�zy��A��5AF�A�4��@��L4�R��A��@�p�. R�Q�R-PPf��@�� ��Ah���=H�9=Ƨ�=�^5=�>P��>���=��,d_�,P�� ���C��<(�U\� 4����_[����A@��?�� pO�_xM�_o0o�ȡT <ofo ovo�o~o�o�o�|I>��y�b��R=���=��yzq���G�G��� � ��!�!�N�Ut@�T��V���uB�� B��B��B%�!����~'���u����q�q6|�\@�&���g���)PB3p�B�B A�@�p"���m���<���  ��e<��)N�3���?���6_�67<�U6[�����C�	��	(@B���]�l���r�ݏ�ȏ��x�"������C3��9 O��C2��@C����q�쏕��������ݟȟN�PB>��)'<�ٗ�����ܿ�*xM��=���CT_CONFIG K�>m�eg7Ų��STBF_TTS��
YɈ�Ȱ��������MAU��N����MSW_CF\�L��  ���OCV7IEW��M�������A�S�e�w��� ����/�Ŀֿ���� ϭ�B�T�f�xϊϜ� +�����������,� ��P�b�t߆ߘߪ�9� ��������(��L� ^�p�����G��� �� ��$�6���Z�l�`~�������D�RC�	N(E��!P�����!�E4iX���S�BL_FAULT� O����GP�MSK���P�TD?IAG P`��q�o��o�U�D1: 6789?012345t�n���P*�Sew �������/ /+/=/O/a/s/2����R
B�/�TR'ECP�
? )�+A>?P?b?t?�? �?�?�?�?�?�?OO (O:OLO^O�/�/�/�O��UMP_OPT�ION����ATR�袒��	�EPME����OY_TEMP�  È�3B��5P��TUN�I͠��5QܦYN_?BRK Q��?EDITOR�A�A�_�R_� ENT �1R��  ,�&PROG A?NIE2 M�Q�_:�D�PICK�_o� &DROP��_3o`
ZEROW#o`o&}�os��to�o�o�o�o�o �o/SeL� p�������  �=�$�a�H�p���~� ����ߏ�؏����P�MGDI_STA�HU$�5Q}UNC;�1S� �dO��v�
�N
�Nd�Oݟ�� �%�7�I�[�m���� ����ǯٯ����!� 3�E�W��En������� ��ʑ��ؿ���� � 2�D�V�h�zόϞϰ� ��������
��.�@� ��g�q߃ߕߧ����� ������%�7�I�[� m����������� ���!�3�E�_�i�{� �������������� /ASew�� �����+ =W�Es����� ���//'/9/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?Oak? }?�?E?��?�?�?�? OO1OCOUOgOyO�O �O�O�O�O�O�O	__ -_G?Y?c_u_�_�_�? �_�_�_�_oo)o;o Mo_oqo�o�o�o�o�o �o�o%7Q_[ m��_���� ��!�3�E�W�i�{� ������ÏՏ���� �/�IS�e�w���� ����џ�����+� =�O�a�s��������� ͯ߯���'�A�3� ]�o���������ɿۿ ����#�5�G�Y�k� }Ϗϡϳ��������� ��9�K�U�g�yߋ� ������������	�� -�?�Q�c�u���� ������������C� M�_�q����ߧ����� ����%7I[ m������ �!;�EWi{ ��������/ ///A/S/e/w/�/�/ �/�/�/�/�/??3 !?O?a?s?��?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_+?=?G_Y_k_ !_�?�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	#_ 5_?Qcu�_�� ������)�;� M�_�q���������ˏ ݏ���-7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� %�/�A�S�e��q��� ����ѿ�����+� =�O�a�sυϗϩϻ� ���������9�K� ]�w����ߥ߷����� �����#�5�G�Y�k� }������������ �'�1�C�U�g��ߋ� ������������	 -?Qcu��� ����m��); M_y������ ��//%/7/I/[/ m//�/�/�/�/�/�/ �/!?3?E?W?q{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O?�O+_ =_O_i?__�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o__#5G�os_ }������� ��1�C�U�g�y��� ������ӏ��o� -�?�Q�ku������� ��ϟ����)�;� M�_�q���������˯ ݯ�	��%�7�I�c� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ��������� �/�A�[�M�w߉ߛ� �߿���������+� =�O�a�s����� ���������'�9�S� e�o������������� ����#5GYk }�������� 1C]�gy� ������	// -/?/Q/c/u/�/�/�/ �/�/I�??)?;? U_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�/ �O_!_3_M?W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�O�o+ E_;as���� �����'�9�K� ]�o���������ɏ�o� �$ENETM�ODE 1TFu��  
�`�`�e�"���RROR_PRO/G %��%�fe��r�@�TABLE  ��P��ß՟��@�SEV_NU�M �  ��	��@�_AU�TO_ENB  q,��=�_NO�� U��!���  *�]��]��]��]��+\�v���<��6�FLTR"�4��HIS��a�/�_�ALM 1V��� ��d]��`+ ��6�H�Z�l�~������_��<�  ���[�"�պ�TCP_�VER !��!�]���$EXTLO�G_REQ֦�-�'�SIZ0�"�SkTKM�K��$¿TOL  �aD�zޢ�A "�_BWD��������'�v��DI�� WFu��� ��a��S�TEP�������O�P_DOo���FD�R_GRP 1X����d 	пm�"��^�n&����c?��$,�MT� ��$ �����^ӳ����^�B�8 B���!C ��B��"dB\�vB%���� $B`��B���Aб�A�e(A�������:�%�^�I���m���  A,��fAt�>(������`
 M��	����ⲉ� ������?�*�c����A@����@�33K@�������@����L�����^�F@ ��E��������L�FZ!D��`�D�� BT��@������?�  M��6����u��5�?Zf5�ES�����e�����J� 9���`�Z�yw�>x�F�EATURE �YFu��&��LR Handl�ingTool ���bEngl�ish Dict�ionary�4�D St� ard���Analog� I/O#,gle Shift?�uto Soft�ware Upd�atedmati�c Backup��	�ground� Edit� �C_amera:F>�Common calib UI���n��Moni�tor�tr� R�eliabS�D�HCP��
Dat�a Acquis��%)iagnos��7?+ocume�nt Viewe�"''ual Ch�eck Safe�ty��hanc�ed��
�%s� F�r��xt. D7IO �fiu$�'wend� Err QLt"	=�'s9r5��  ���
FCTN_ Menu� v##�[7TP InJ0f�acq5�GigE��>�5�p Mas_k Exc� g�'�HT�0Proxy� Sv�$�6igh�-Spe� Ski��6m � mmun�ic�onsHu�rh0J0:/;�2connect 2:H�ncr�0struH8Ja@e�!� Jt%��KAREL C�md. L�0ua��8�CRun-Ti�� Env�HK0el� +�s�S/W��License��#�,0Book(System)�
MACROs,�2?/OffseZUaH� w8/"PMR D�s.M}M@!l�,�MechStop"�1tQ@Y"Ui2V©Vx� 7�L^od>Twitch�_aS�h!.BV�[Optm�oaS�0fi�^aVg�0GUulti-T��0��	PCM f�unkG�ia�Pti�z~h�goV$RegeiPr@�fri� �F�k�f8Num �Sel�U�i�  Adju@�n qV1}tatu�aI�*��RDM Robo}tscove�ueav`� Fre�q AnlyGRem�P�!n�u�rServo� �P�?SNPX b�B[;SN�0Cli�!�WLibr(�� Q �T:��vo�@th0�ssag~e�� 0l5Q&�/I�=���MILIB����P� Firmu��P�h3Acc��TPsTX4/��eln5P�Ǐ���1U��orq}uTimula!4�E�u�PPa�A���!!c&�0ev.́�mri� �USR EVNTğ�֐nexcept�� �pn�#ѕ�(@VEC�rBB�XVU �6��G�:�A�S�S9C�y�SGE�����UI&Web Pl`vǮ�q0O��0�$��!?6ZDT Ap�plD�
iP0a|!�:� Grid�qplay=����W�R-�.��h!N��B<^P}200iV4+�scii�1rLosad� �Upl��8�f@I�Pat�V�ycS�B�`��� \6�RL��� ۩�5MIo Dev�@ (�q�R�f�?�gsswo�!�_64MB �DRAMM���FR9O�Ͼell:�#sh��#�c.k ղrp��5�tySs
r7̬r'`.?+�p�!X"=-o� 2�a5port�.�p�r q�-T1 �{]P���No m�pc�$筴OL��Sup���Fa�hOPC-UA�l�T �2eϓ�9S0�0croa|�s�:����~���ues�t�uS��e2te�xV��up�1�#��P�P�00�oVirt��!�sR�stdpn�Û�� SWIMEoST f F0��������������� �� MDVp z������ 
I@Rlv� �����/// E/</N/h/r/�/�/�/ �/�/�/???A?8? J?d?n?�?�?�?�?�? �?O�?O=O4OFO`O jO�O�O�O�O�O�O_ �O_9_0_B_\_f_�_ �_�_�_�_�_�_�_o 5o,o>oXobo�o�o�o �o�o�o�o�o1( :T^����� ��� �-�$�6�P� Z���~�������Ə� ���)� �2�L�V��� z����������� %��.�H�R��v��� ����������!�� *�D�N�{�r������� ���޿���&�@� J�w�nπϭϤ϶��� ������"�<�F�s� j�|ߩߠ߲������� ���8�B�o�f�x� ������������ �4�>�k�b�t����� ��������0 :g^p���� ��	 ,6c Zl������ /�/(/2/_/V/h/ �/�/�/�/�/�/?�/ 
?$?.?[?R?d?�?�? �?�?�?�?�?�?O O *OWONO`O�O�O�O�O �O�O�O�O__&_S_ J_\_�_�_�_�_�_�_ �_�_�_o"oOoFoXo �o|o�o�o�o�o�o�o �oKBT�x �������� �G�>�P�}�t����� ����������C� :�L�y�p��������� �ܟ���?�6�H� u�l�~��������د ���;�2�D�q�h� z�������ݿԿ� � 
�7�.�@�m�d�vϣ� �Ϭ����������3� *�<�i�`�rߟߖߨ� ���������/�&�8� e�\�n�������� ������+�"�4�a�X� j��������������� ��'0]Tf� �������# ,YPb��� �����//(/ U/L/^/�/�/�/�/�/ �/�/�/??$?Q?H? Z?�?~?�?�?�?�?�? �?OO OMODOVO�O zO�O�O�O�O�O�O_ 
__I_@_R__v_�_ �_�_�_�_�_ooo Eo<oNo{oro�o�o�o �o�o�oA8 Jwn����� ����=�4�F�s��j�|�����̍  H551��z�2�R782�{50�J614��ATUP�545z�6�VCAM�oCUIF�28H��NRE�52;�R�63�SCH�DwOCV��CSU��869�0�EI�OCl�4��R69�;�ESET$�:�J�7:�R68�MA{SK�PRXYT�]7�OCO�3$�h�����37�J6
��53��He�LCH^�OPLG$�0O��MHCR �S��M�ATk�MCS#�0���55�MDSW��B�OPB�MPR�C���s�0�PCM�S�5J������s�5�1/�51{�0/�P�RS�697�FR�DG�FREQ�M�CN�93�SN�BAx�f�SHLB��M
ǀ���2�H{TC#�TMIL�TPA˖TPT�X<�EL۶����8������J95_�T�UTC�UEV�U�EC�UFRG�V�CC��OǦVIP�G�CSCk�CSGtk���I�WEB#�7HTT#�R6v����CG6�IG�IP�GS\�RCG�DGnB�H75/�R7�]Ry�R66O�2O��R6�R55��4���5��D06�F��CLI3�.�CMqS˖0�#�STY�ǋTO7�7��t�_�O�RSǦ��M��NOM˖OL�$����OPIs�SEND��L��Sy�ETS�sּ�S�CPk�FV�R˖IPNG�Gene�È6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�P�b�t��������� ������(:L�^p�����	�  H55�1��2�
R78�2�50�	J61�4�	ATUP5�456�	VCA�M�	CUIF2�8lNRE�
52�[R63�SCH��	DOCV�CS]U�
8690+�EIOC�4R{69[ESET<vZJ7ZR68�
�MASK�	PRXuY|7�
OCOL,�3<X 3�*J�653�H�,L{CH�*OPLG<�0�*MHCR�*S�J;MAT�MCS�;0[+55+MD�SW�;�+OP�+M�PR�*��,0PCM{5KX +X0��+51K51[L0nKPRSK+69�*�FRDkFREQn�
MCN�
93�SNBA��+SH�LB�JM[��<2�HTC;TMI�L��TPA*T7PTX\ZEL�JX0��8
�
J95�TUT�*UEV�K*UEC�*UFR�kVCC+lOk:V�IPkZCSC�ZC�SG��I�	WE�B;HTT;R6l��\CG�kIG�koIPGS�jRCkZ�DG�+H75KRu7:+RYLR66�,�2�*R6�R55�k|4�[5�{D06:+F�|CLI�<J�CMS*�p;ST-Y[kTO�k7����ORSk:x Mn�LNOM*OL�;��0�OPI�jSE�ND�
L:kSY�EcTS�j {[CP�wFVR*IPNkZGene��R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt������� �STD�LANG��	' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__�)_;_M___q_�ZRB=T�OPTN�_�_��_�_�_DPN �oo*o<oNo`oro �o�o�o�o�o�o�o~ted � �>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�X�j� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FXj |�������p��0�B�  �K��i�{�������Í9�9ʅ�$FEAT�_ADD ?	��������  	ǈ��,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n��������������� ��"4FXj| ������� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�DEMO Y��?   ǈ1] '_9_f_]_o_�_�_�_ �_�_�_�_�_,o#o5o boYoko�o�o�o�o�o �o�o�o(1^U g������� �$��-�Z�Q�c��� ����Ə��Ϗ�� � �)�V�M�_������� ��˟����%� R�I�[���������� ǯ����!�N�E� W���{�������ÿݿ ����J�A�Sπ� wω϶ϭϿ������ ��F�=�O�|�s߅� �ߩ߻�������� B�9�K�x�o���� ����������>�5� G�t�k�}��������� ����:1Cp gy�����  �	6-?lcu �������/ 2/)/;/h/_/q/�/�/ �/�/�/�/�/?.?%? 7?d?[?m?�?�?�?�? �?�?�?�?*O!O3O`O WOiO�O�O�O�O�O�O �O�O&__/_\_S_e_ �_�_�_�_�_�_�_�_ "oo+oXoOoao�o�o �o�o�o�o�o�o 'TK]���� ������#�P� G�Y���}��������� ׏����L�C�U� ��y�������ܟӟ� �	��H�?�Q�~�u� ������دϯ��� �D�;�M�z�q����� ��Կ˿ݿ
���@� 7�I�v�m�ϙϣ��� ��������<�3�E� r�i�{ߕߟ������� ����8�/�A�n�e� w������������ �4�+�=�j�a�s��� ������������0 '9f]o��� �����,#5 bYk����� ���(//1/^/U/ g/�/�/�/�/�/�/�/ �/$??-?Z?Q?c?}? �?�?�?�?�?�?�? O O)OVOMO_OyO�O�O �O�O�O�O�O__%_ R_I_[_u__�_�_�_ �_�_�_oo!oNoEo Woqo{o�o�o�o�o�o �oJASm w������� ��F�=�O�i�s��� ����֏͏ߏ��� B�9�K�e�o������� ҟɟ۟����>�5� G�a�k�������ίů ׯ����:�1�C�]� g�������ʿ��ӿ � ��	�6�-�?�Y�cϐ� �ϙ��Ͻ�������� 2�)�;�U�_ߌ߃ߕ� �߹��������.�%� 7�Q�[������ ��������*�!�3�M� W���{����������� ����&/IS� w������� "+EO|s� ������// '/A/K/x/o/�/�/�/ �/�/�/�/??#?=? G?t?k?}?�?�?�?�? �?�?OOO9OCOpO gOyO�O�O�O�O�O�O _	__5_?_l_c_u_ �_�_�_�_�_�_oo o1o;oho_oqo�o�o �o�o�o�o
- 7d[m���� �����)�3�`� W�i�������̏ÏՏ ����%�/�\�S�e� ������ȟ��џ���� �!�+�X�O�a����� ��į��ͯ����� '�T�K�]��������� ��ɿ������#�P� G�Yφ�}Ϗϼϳ���������   �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�O�O �O__/_A_S_e_w_ �_�_�_�_�_�_�_o o+o=oOoaoso�o�o �o�o�o�o�o' 9K]o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ����/�A�S�e�w� ������������ �+�=�O�a�s����� ����������' 9K]o���� ����#5G Yk}����� ��//1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O��O�O�O�O_Y  XQ/_A_S_ e_w_�_�_�_�_�_�_ �_oo+o=oOoaoso �o�o�o�o�o�o�o '9K]o�� �������#� 5�G�Y�k�}������� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���������ϯ�� ��)�;�M�_�q��� ������˿ݿ��� %�7�I�[�m�ϑϣ� �����������!�3� E�W�i�{ߍߟ߱��� ��������/�A�S� e�w��������� ����+�=�O�a�s� �������������� '9K]o�� ������# 5GYk}��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{��������� ������/AS ew������ �+=Oas �������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? 5?G?Y?k?}?�?�?�? �?�?�?�?OO1OCO UOgOyO�O�O�O�O�OP�O�O	_QPX 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o��� ������ɏۏ���� #�5�G�Y�k�}����� ��şן�����1� C�U�g�y��������� ӯ���	��-�?�Q� c�u���������Ͽ� ���)�;�M�_�q� �ϕϧϹ�������� �%�7�I�[�m�ߑ� �ߵ����������!� 3�E�W�i�{���� ����������/�A� S�e�w����������� ����+=Oa s������� '9K]o� �������/ #/5/G/Y/k/}/�/�/ �/�/�/�/�/??1? C?U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o �o�o�o�o�o�o! 3EWi{��� ������/�A� S�e�w���������я �����+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ���� #�5�G�Y�k�}����� ��ſ׿�����1� C�U�g�yϋϝϯ����������	���$F�EAT_DEMO�IN   Ԁ�K�� �3�IND�EX@�Oш3�I�LECOMP �Z������N�.�w�SETU�P2 [��~���  N ���t�_AP2BCK� 1\��  #�)�����%��� ����H����t� ��'����]���� �(���L���p���� ��5�����k� ��$ ��1Z��~�� C�g��2� Vh���?� �u
/�./@/�d/ ��/�/)/�/M/�/�/ �/?�/<?�/I?r?? �?%?�?�?[?�??O &O�?JO�?nO�OO�O 3O�OWO�O�O�O"_�O F_X_�O|__�_�_A_ �_e_�_o�_0o�_To �_ao�oo�o=o�o�o so�o,>�ob�o ��'�K�o�������P�� 2>��*.VR�g��p*j����s������uQ�PC��pOFR6:֏���;�ʋT_�_�q� �\����B�,����v*.FT���q	�������C�қSTM @c�l�w��d����p�iPendant Panel��қH������该�3�L�ӚGIFV������l�)�;�пӚJPG ڿϋ�𿭿��T�ˊ#JS^χ��p�u��2�%
JavaS�cript��޿C�S��ߊ��ϵ� %�Cascadi�ng Style Sheets7���p
ARGNAMOE.DTf��|���\z�8ߚ��Ի�g�>��DISP*�ߔ߀����>���0�?���	?PANEL15��%�����ﵯǯu�2����������o�z�3;������L�^���z�4��%�������wr�TPEIN�S.XML~�:�\�PbCust�om Toolb�ar���PASS�WORDC�~F�RS:\� %�Passwor�d ConfigW��4�/�ԝ[ U�/qֱ䘯���/��b_/v���/%@J(�/g/y/?'2T/ =?H(+?�/�/�?��?��/U5�?o?�?O'3 \?EOH(3O�?O�O�� �O�?]E�OwO�O_'4dOM_H(;_�O_�_ �_�OeU�__�_&o �Jo�no���o3o �oWo�o�o�o"�oF X�o|��A� e���0��T�� M������=�ҏ�s� ���,�>�͏b�񏆟 �'���K���o�ٟ� ��:�ɟ^�p�����#� ��ʯY��}������ H�ׯl���e���1�ƿ U������ ϯ�D�V� �z�	Ϟ�-�?���c� �χ���.߽�R���v� ��߬�;�����q�� ��*����`��߄�� }��I���m����� 8���\�n����!��� E�W���{���	F ��j����/�S ����B�� x�+��a��,�$FILE_�DGBCK 1\������� < �)�
SUMMARY�.DG/�]MD:�:/z/�Dia�g Summar�y{/([CONSLOGp/S/e!�/�/�!�Console� log�/�\TPOACCN�/Y?%A?�~?�%TP Accountin ?��Y@6:IPKD?MP.ZIP�?��
�?O�%�0Exc?eptionO�#*�_\O�bQJO��_1FR DT Files�O�<f �MEMCHECK�t?�/i/_1Me�mory Dat�a_�l�)	FTP�/f_�Oj_�W1mme`T�BD�_�L >I�)ETHERNET�_��A�_o�!�Etherne�t 0figur�a&O�}QDCSV�RF�_m__�oQ�%]` veri?fy all�o��M.cXeDIF�F�ovo�o P%=�hdiff�g|�A]`CHG01��o��a5��b- `y2��&�1��gr3������ <�я`�V�TRNDIAG.�LS֏����.�!Q�� Ope>c L�og �!nost�icCW��)oVDEV�DA}O������aVis~Q�DeviceX�e�IMG��?�����4�7�ʔImag�֟c�UP{�ES�z��FRS:\�z��O@Updates List����"�FLEXEVENo�%�>��a�� UIF E�v�QU�?�  ,��sz)
PSRB?WLD.CMj���������0PS_ROBOWEL�_��*�HADOW�4��+�D�SSh�adow Chasng�ODVa��?RCMERR<�!��3���S��CFG� ErrorАt�ailk� a���B��SGLIB��ϧϹ�N�!Q� �St?`_�����):�ZDU_��7����WZDT�ad�n����NOTI�bo�߽�R�UNotific?b��t���AGXbGIGE���/�A���]�Gig�EZ�d��N�A� �-��Q��^���� ��:�����p���) ;��_����$� H�l��7� [m�� ��V �z/!/�E/�i/ �v/�/./�/R/�/�/ �/?�/A?S?�/w?? �?�?<?�?`?�?�?O +O�?OO�?sO�OO�O 8O�O�OnO_�O'_9_ �O]_�O�__�_�_F_ �_j_�_o�_5o�_Yo ko�_�oo�o�oTo�o xo�oC�og�o ��,�P��� ��?�Q��u���� (���Ϗ^�󏂏�)� ��M�܏q������6� ˟ݟl����%���2� [��������D�ٯ h������3�¯W�i� �������@����v� Ϛ�/�A�пe����� ��*Ͽ�N����τ�� ��=���J�s�ߗ�&� ����\��߀��'�� K���o����4��� X������#���G�Y� ��}������B���f� ����1��U��b ��>��t	��$FILE_�FRSPRT  ���� ����$MDO?NLY 1\8� ? 
 ��{ �������� ///�S/�w/�// �/</�/�/r/?�/+? �/8?a?�/�??�?�? J?�?n?OO�?9O�? ]OoO�?�O"O�OFO�O �O|O_�O5_G_�Ok_ �O�_�_0_�_T_�_�_ �_o�_Co�_Poyo"?VISBCKV@>e*.VD�o�o�8`FR:\�`I�ON\DATA\��oZb8`Vis�ion VD file�oo>Pfo t^o�'��]� ��(��L��p�� ���5�ʏ܏�� ��� $���5�Z��~���� ��C�؟g�������2� ��V�h�#������?� ���u�
���.�@�ϯ�d�󯈿�)���L�UI_CONFIoG ]8�a>ɻ $ ��[{8 �2�D�V�h�z����|x�������� ����
ܠ�-�?�Q�c� u�߆߽߫������� ���)�;�M�_�q�� ������������ %�7�I�[�m������ ����������!3 EWi ���� ��~/AS e������h �//+/=/O/�s/ �/�/�/�/�/d/�/? ?'?9?K?�/o?�?�? �?�?�?`?�?�?O#O 5OGO�?kO}O�O�O�O �O\O�O�O__1_C_ �Og_y_�_�_�_�_X_ �_�_	oo-o�_>oco uo�o�o�oBo�o�o�o )�oM_q� ��>����� %��I�[�m������ :�Ǐُ����!��� E�W�i�{�����6�ß ՟�������A�S� e�w��� �����ѯ� �����+�=�O�a�s� �������Ϳ߿�� ��'�9�K�]�oρ�� �Ϸ��������ϖ�#� 5�G�Y�k�}�ߡ߳� �������ߎ��1�C�PU�g�y�	���x������$FLUI_�DATA ^���������RESUL�T 2_����� �T�/w�izard/gu�ided/ste�ps/Expert��"�4�F�X�j�|����������������Continue with G��ance��1C Ugy������ ��-����0 ����l��$���ps� o������� �/#/5/���\/n/ �/�/�/�/�/�/�/�/ ?"?4?F>$(:Jrip�X�? �?�?�?OO*O<ONO `OrO�OC/�O�O�O�O �O__&_8_J_\_n_��_�_Q?c?�_�?E�J�TimeUS/DST�_"o4oFo Xojo|o�o�o�o�o�o~��Enabl 
.@Rdv���������� �_��_�_f24 or���������̏ޏ ����&��o�o\�n� ��������ȟڟ��� �"�4����)�;�M�zon
`7�ʯܯ � ��$�6�H�Z�l��~���EST E�a�rn Stand������ӿ��� 	��-�?�Q�c�uχ�� ��t�f�x��:���acces �?�+�=�O�a�s߅ߠ�ߩ߻�������n�ect to N?etwork��� %�7�I�[�m����P������ȘA���Ⱥ��ϊ�!��`In�troduction��t��������� ������(�OL ^p������ � $5�_��P*����VEditor5����
/�/./@/R/d/v/5 �Touch Pa�nel � (recommen�P)�/�/�/�/�/?#?@5?G?Y?k?}?�̬P� ^�?�B�?OO/O AOSOeOwO�O�O�O�O �O<�O__+_=_O_ a_s_�_�_�_�_�_�Y�0�?�:�?o�? EoWoio{o�o�o�o�o �o�o�o�OAS ew������ ���+��_�_op� 2o������͏ߏ�� �'�9�K�]�o�.�� ����ɟ۟����#� 5�G�Y�k�}�<���`� ¯�������1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ��ώ��� ���֯;�M�_�q߃� �ߧ߹��������� %��I�[�m���� �����������!��� B��f�(�*������� ������/AS ew6����� �+=Oas 2��V�����/ /'/9/K/]/o/�/�/ �/�/�/��/�/?#? 5?G?Y?k?}?�?�?�? �?����?O�CO UOgOyO�O�O�O�O�O �O�O	__�/?_Q_c_ u_�_�_�_�_�_�_�_ oo�? O�?Dono0O �o�o�o�o�o�o %7I[m,_�� ������!�3� E�W�i�(o:oLo^o�� �o�����/�A�S� e�w���������~� ����+�=�O�a�s� ��������ͯ������ �ԏ9�K�]�o����� ����ɿۿ����П 5�G�Y�k�}Ϗϡϳ� ����������ޯ� �d�&��ߝ߯����� ����	��-�?�Q�c� "�t���������� ��)�;�M�_�q�0� ��T߶�x����� %7I[m�� ������!3 EWi{���� �����/��//A/S/ e/w/�/�/�/�/�/�/ �/??�=?O?a?s? �?�?�?�?�?�?�?O O�6O�ZO/O�O �O�O�O�O�O�O_#_ 5_G_Y_k_*?�_�_�_ �_�_�_�_oo1oCo Uogo&O�oJO�o�o�_ �o�o	-?Qc u����|_�� ��)�;�M�_�q��� ������xo�o�o�� �o7�I�[�m������ ��ǟٟ�����3� E�W�i�{�������ï կ����ʏ��8� b�$���������ѿ� ����+�=�O�a� � �ϗϩϻ�������� �'�9�K�]��.�@� R���v��������#� 5�G�Y�k�}���� r���������1�C� U�g�y����������� �ߤ���-?Qc u������� ��);M_q� ������// ������X//�/�/ �/�/�/�/�/?!?3? E?W?h?�?�?�?�? �?�?�?OO/OAOSO eO$/�OH/�Ol/�O�O �O__+_=_O_a_s_ �_�_�_�_�O�_�_o o'o9oKo]ooo�o�o �o�ovO�o�O�o�O# 5GYk}��� ������_1�C� U�g�y���������ӏ ���	��o*��oN� ���������ϟ�� ��)�;�M�_���� ������˯ݯ��� %�7�I�[��|�>��� ��v�ٿ����!�3� E�W�i�{ύϟϱ�p� ��������/�A�S� e�w߉ߛ߭�l����� ���ƿ+�=�O�a�s� ������������ ��'�9�K�]�o����� ��������������� ��,V�}��� ����1C U�y����� ��	//-/?/Q/ "4F�/j�/�/�/ ??)?;?M?_?q?�? �?�?f�?�?�?OO %O7OIO[OmOO�O�O �Ot/�/�/�O�/!_3_ E_W_i_{_�_�_�_�_ �_�_�_�?o/oAoSo eowo�o�o�o�o�o�o �o�O�O�OL_s �������� �'�9�K�
o\����� ����ɏۏ����#� 5�G�Y�z�<��` şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u�������j�̿��� ���)�;�M�_�qσ� �ϧϹ���������� %�7�I�[�m�ߑߣ� ���������߼��� B���{������ ��������/�A�S� �w������������� ��+=O�p 2��j���� '9K]o�� �d�����/#/ 5/G/Y/k/}/�/�/` ���/�/�?1?C? U?g?y?�?�?�?�?�? �?�?�O-O?OQOcO uO�O�O�O�O�O�O�O �/�/�/ _J_?q_�_ �_�_�_�_�_�_oo %o7oIoOmoo�o�o �o�o�o�o�o!3 E__(_:_�^_� �����/�A�S� e�w�����Zo��я� ����+�=�O�a�s� ������hz� �'�9�K�]�o����� ����ɯۯ���#� 5�G�Y�k�}������� ſ׿�����̟ޟ@� �g�yϋϝϯ����� ����	��-�?���P� u߇ߙ߽߫������� ��)�;�M��n�0� ��TϹ��������� %�7�I�[�m������ ����������!3 EWi{��^�� �����/AS ew������ ���/+/=/O/a/s/ �/�/�/�/�/�/�/� ?�6?��/o?�?�? �?�?�?�?�?�?O#O 5OGO/kO}O�O�O�O �O�O�O�O__1_C_ ?d_&?�_�_^O�_�_ �_�_	oo-o?oQoco uo�o�oXO�o�o�o�o );M_q� �T_�_x_���_� %�7�I�[�m������ ��Ǐُ돪o�!�3� E�W�i�{�������ß ՟矦���>� � e�w���������ѯ� ����+�=���a�s� ��������Ϳ߿�� �'�9���
��.��� R������������#� 5�G�Y�k�}ߏ�N��� ����������1�C� U�g�y���\�nπ� ���	��-�?�Q�c� u��������������� );M_q� ���������� ��4��[m�� �����/!/3/ ��D/i/{/�/�/�/�/ �/�/�/??/?A?  b?$�?H�?�?�?�? �?OO+O=OOOaOsO �O�O�?�O�O�O�O_ _'_9_K_]_o_�_�_ R?�_v?�_�?�_o#o 5oGoYoko}o�o�o�o �o�o�o�O1C Ugy����� ��_��_*��_�c� u���������Ϗ�� ��)�;��o_�q��� ������˟ݟ��� %�7��X��|���R� ��ǯٯ����!�3� E�W�i�{���L���ÿ տ�����/�A�S� e�wω�H���l����� ����+�=�O�a�s� �ߗߩ߻����ߞ�� �'�9�K�]�o��� ���������Ͼ�� 2���Y�k�}������� ��������1�� Ugy����� ��	-����� "��F������ //)/;/M/_/q/�/ B�/�/�/�/�/?? %?7?I?[?m??�?P bt�?��?O!O3O EOWOiO{O�O�O�O�O �O�/�O__/_A_S_ e_w_�_�_�_�_�_�_ �?�?�?(o�?Ooaoso �o�o�o�o�o�o�o '�O8]o�� �������#� 5��_V�oz�<o���� ŏ׏�����1�C� U�g�y���������ӟ ���	��-�?�Q�c� u���F���j�̯��� ��)�;�M�_�q��� ������˿ݿ���� %�7�I�[�m�ϑϣ� �����Ϙ��ϼ��� ��W�i�{ߍߟ߱��� ��������/��S� e�w��������� ����+���L��p� ��F���������� '9K]o�@� ������# 5GYk}<���`� �����//1/C/ U/g/y/�/�/�/�/�/ ��/	??-???Q?c? u?�?�?�?�?�?�� ��?&O�MO_OqO�O �O�O�O�O�O�O__ %_�/I_[_m__�_�_ �_�_�_�_�_o!o�? �?OOxo:O�o�o�o �o�o�o/AS ew6_����� ���+�=�O�a�s� ��DoVohoʏ�o�� �'�9�K�]�o����� ����ɟ�����#� 5�G�Y�k�}������� ůׯ�������ޏC� U�g�y���������ӿ ���	��ڟ,�Q�c� uχϙϫϽ������� ��)��J��n�0� �ߧ߹��������� %�7�I�[�m��ߣ� �����������!�3� E�W�i�{�:ߜ�^��� ������/AS ew������� �+=Oas ���������� /���K/]/o/�/�/ �/�/�/�/�/�/?#? �G?Y?k?}?�?�?�? �?�?�?�?OO�@O /dOvO:?�O�O�O�O �O�O	__-_?_Q_c_ u_4?�_�_�_�_�_�_ oo)o;oMo_oqo0O zOTO�o�o�O�o %7I[m�� ���_���!�3� E�W�i�{�������Ï �o�o�o����oA�S� e�w���������џ� �����=�O�a�s� ��������ͯ߯�� �ԏ���
�l�.��� ����ɿۿ����#� 5�G�Y�k�*��ϡϳ� ����������1�C� U�g�y�8�J�\��߀� ����	��-�?�Q�c� u�����|����� ��)�;�M�_�q��� ���������ߜ߮� ��7I[m�� �������  EWi{���� ���//��>/  b/$�/�/�/�/�/�/ �/??+?=?O?a?s? �/�?�?�?�?�?�?O O'O9OKO]OoO./�O R/�Ov/�O�O�O_#_ 5_G_Y_k_}_�_�_�_ �_�?�_�_oo1oCo Uogoyo�o�o�o�o�O �o�O�O�o?Qc u������� ���_;�M�_�q��� ������ˏݏ��� �o4��oX�j�.����� ��ǟٟ����!�3� E�W�i�(�������ï կ�����/�A�S� e�$�n�H�����~�� ����+�=�O�a�s� �ϗϩϻ�z������ �'�9�K�]�o߁ߓ� �߷�v��������п 5�G�Y�k�}���� �����������1�C� U�g�y����������� ����	��������` "������� );M_�� ������// %/7/I/[/m/,>P �/t�/�/�/?!?3? E?W?i?{?�?�?�?p �?�?�?OO/OAOSO eOwO�O�O�O�O~/�/ �/_�/+_=_O_a_s_ �_�_�_�_�_�_�_o �?o9oKo]ooo�o�o �o�o�o�o�o�o�O 2�OV_}��� ������1�C� U�g�x��������ӏ ���	��-�?�Q�c� "��F��jϟ�� ��)�;�M�_�q��� ������x�ݯ��� %�7�I�[�m������ ��t�ֿ��������3� E�W�i�{ύϟϱ��� �������ʯ/�A�S� e�w߉ߛ߭߿����� ���ƿ(��L�^�"� ������������ �'�9�K�]�߁��� ������������# 5GY�b�<�� r����1C Ugy���n�� ��	//-/?/Q/c/ u/�/�/�/j���/ ?�)?;?M?_?q?�? �?�?�?�?�?�?O� %O7OIO[OmOO�O�O �O�O�O�O�O�/�/�/ �/T_?{_�_�_�_�_ �_�_�_oo/oAoSo Owo�o�o�o�o�o�o �o+=Oa _ 2_D_�h_���� �'�9�K�]�o����� ��doɏۏ����#� 5�G�Y�k�}������� r������1�C� U�g�y���������ӯ ������-�?�Q�c� u���������Ͽ�� �ğ&��J��qσ� �ϧϹ��������� %�7�I�[�l�ߑߣ� �����������!�3� E�W��x�:Ϝ�^��� ��������/�A�S� e�w�������l����� ��+=Oas ���h������� �'9K]o�� ��������#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/�?�@? R?/y?�?�?�?�?�? �?�?	OO-O?OQO/ uO�O�O�O�O�O�O�O __)_;_M_?V?0? z_�_f?�_�_�_oo %o7oIo[omoo�o�o bO�o�o�o�o!3 EWi{��^_�_ �_���_�/�A�S� e�w���������я� ���o�+�=�O�a�s� ��������͟ߟ� ���H�
�o����� ����ɯۯ����#� 5�G��k�}������� ſ׿�����1�C� U��&�8���\����� ����	��-�?�Q�c� u߇ߙ�X��������� ��)�;�M�_�q�� ���f�xϊ����� %�7�I�[�m������ ������������!3 EWi{���� �������> � ew������ �//+/=/O/`s/ �/�/�/�/�/�/�/? ?'?9?K?
l?.�? R�?�?�?�?�?O#O 5OGOYOkO}O�O�O`/ �O�O�O�O__1_C_ U_g_y_�_�_\?�_�? �_�?�_o-o?oQoco uo�o�o�o�o�o�o�o �O);M_q� �������_� �_4�F�
m������ ��Ǐُ����!�3� E�i�{�������ß ՟�����/�A� � J�$�n���Z���ѯ� ����+�=�O�a�s� ����V���Ϳ߿�� �'�9�K�]�oρϓ� R���v����Ϭ��#� 5�G�Y�k�}ߏߡ߳� �����ߨ���1�C� U�g�y�������� ��϶�����<���c� u��������������� );��_q� ������ %7I��,��P� �����/!/3/ E/W/i/{/�/L�/�/ �/�/�/??/?A?S? e?w?�?�?Zl~�? �OO+O=OOOaOsO �O�O�O�O�O�O�/�O _'_9_K_]_o_�_�_ �_�_�_�_�_�?o�? 2o�?Yoko}o�o�o�o �o�o�o�o1C Togy����� ��	��-�?��_`� "o��Fo����Ϗ�� ��)�;�M�_�q��� ��T��˟ݟ��� %�7�I�[�m����P� ��t�֯�����!�3� E�W�i�{�������ÿ տ翦���/�A�S� e�wωϛϭϿ����� ���Ư(�:���a�s� �ߗߩ߻�������� �'�9���]�o��� ������������#� 5���>��b���N߳� ��������1C Ugy�J��� ��	-?Qc u�F���j����� //)/;/M/_/q/�/ �/�/�/�/�/�?? %?7?I?[?m??�?�? �?�?�?����0O �WOiO{O�O�O�O�O �O�O�O__/_�/S_ e_w_�_�_�_�_�_�_ �_oo+o=o�?O O �oDO�o�o�o�o�o '9K]o�@_ �������#� 5�G�Y�k�}���No`o�roԏ��$FMR�2_GRP 1`���� ��C4  B�.�p	 �p�0���F@ F�E���Q�F���C��L��FZ!D�`��D�� BT���@���^�?� � �����6��������5�Zf�5�ESΑ^�A�3  ���BH��\�~�@�33@��	 ����@�Q���@�g�]�Q����<��z�<�ڔ=�7�<�
;;�*�<��^��8ۧ�9k'V�8��8����7ג	8(�� ~�����=�(�a�L�����w�_CFG a�T0���ӿ�|����NO �/
F0+� 0����RM_CHKTYP  �p	������ROMF�_MsINL��s��x�u�7�X�SSB���b�� ��ϙu�����ϝ��TP_DEF_O/W  �t	��ǟIRCOMK�����$GENOVRD�_DOm��q*�T[HRm� dG�d0�o_ENB� 0ЯRAVC��c���� �>�����v����^����.� ���OU��i��3�.��.�< u�����,�z����sC�  D����l�d�$�@��B�/���1�m��ϑ�SMT���j��������$�HOSTC��1k������� kMC�t�����v  27.0z 1��  e�� BTfx�
0�������	anonymous 4FXj|�r���������)
/ /./@/R/�v/�/�/ �/�i/�/??*? <?N?����?�/�? ��?�?OO�/�?JO \OnO�O�?�O�/�O�O �O�O_S?�Ow?�?j_ �O�?�_�_�_�_�_+O oo0oBoTow_�O�O �o�o�o�o�o'_9_K_ ]__o5�_t��� ��_����(�K }o�op����������o 13�$�gH�Z� l�~������Ɵ؟� ���Q��D�V�h�z� ��Ϗ�󏥯���;� �.�@�R�d������� ������%���*� <�N�`ϣ���ǯ��ۿ �������&�i�J� \�n߀ߒߵ�7�����������"�o���EN�T 1l��� � P!��s�  u�a�������� ��
������?�d�'� ��K���o��������� ��*��Nr5� Yk����� 8�1n]�U� y����/4/� X//|/?/�/c/�/�/��/�/�/?�/B?:?QUICC0O?+?=?�?a41�?{?�?�?�a42�?�?�?>O!?ROUTER?OO�-O�O!PCJO�G�OjO!19�2.168.0.�10h?]3CAMP�RT�O�O!�E1�@_�FRTXO
__�}_C�NAME �!P�!ROBO��O�_S_CFG �1kP� ��Auto-s�tarted��FTP��a�Ϧ� Ao��eowo�o�o�oF� �o�o�o*o�oO as���r��_o o�'Io�<�N�`� r�5������̏ޏ� ���&�8�J�\�n�g� yϋϝ�鏿����� "�4�F�	�j�|����� ��՟W������0� B�������������� ҿ�����ݯ>�P� b�tφϩ�+ϼ����� ����Y�k�}�/ߑ� ��ſ�߸������߱� �$�6�H�k�l��ߐ� ���������-�?�Q� 2�e�V���z������� s�������
?��� ;dv������ �%�9[�<N` r�G����� �&/8/J/\/n/�/ ������//? "?4?F?X?/|?�?�? �?�?�/i?�?OO0O�BOTO�Z_ERR �m�Z\OlFPDU�SIZ  �0^�0��D>�EWR�D ?�U�!� � guest�6�O�O __$_�6_�TSCD_GR�OUP 3n�\ u�Q�9IFT|^w$PA|^OMP|^w |^_SH|^�ED�_ $C|^C�OMn@TTP_A�UTH 1o{K� <!iPen�danBWMn�[�2��q!KAREL�:*MoVohmKC�}o�o�ou`VISION SETfP�o�o�v!,rc P>hb�������~dCTRL Kp{M6��1
1�FFF9E3���$FRS:D�EFAULT[��FANUC W�eb Server[�I��"d�O�D��я�����+�jDW�R_CONFIGw qkU�B�c[�lAIDL_C_PU_PCz��1sB�� �� BH���MIN��sQ��GNR_IOuA�B�0�H���NPT_SIM�_DOӖݛSTAL_SCRNӖ� �ޚTPMOD�NTOL�ݛ��R�TY������` `E�NB�sS��OL_NK 1r{KxP ����ɯۯ������_MASTEҐy��5���SLAVE �s{KH D��S�RAMCACHE�/�A�"aO_CFGq�����UO�`����?CMT_OPz�ՒJǳYCLp���t�_ASG 1t`��A
 �6�H�Z� l�~ϐϢϴ����������� ��	�NUMj�CI
��IPn����RTRY_CN8ҿ���_UP_��A�����E ������]u)�  06������RCA_ACC� 2vk[  R��� C� ��� 4@� W6��026��2� ��#���  z�D���BUF001 2wk[�= Bu��uW0Q��b��q��U��䑖䢖䱖�U�і���������"��1����Wu0*��J@ku0H�_�z���������u0��\@����u0�" S�u0�#�Q����n�0u0Ch1W�An�Pn�an�Upn�n��n��n�~M��f�پ���f`������,u0�rx�D��(gd�u0Pm���u0&@N���N��\p��������������o��  o�R���RU�.�.�.�.-���S�����	�s�2�������������t� x������ ���������� �������������s��$�u ��,��4��=��E��M�t� �T�t� �\�Ye��l� �t�q}�Y��y�� q��q��q��q���q��qM��^����'�M���u0�Z����BH2����1�C8��3HA����	"  	" 	" 	"% &, ��49"= 9"E 9"M �9"U ��\�e s{(lph�t��s�3����"�� ��"�� ����"�� ��"����"���2 ��2�2�2 %�2-�� 5�C2E� S2U�� ]�2e�=� m�JPu�=���JP�� �=���=���=� _4��=�� �� �� �2���2���2���2�� �2#�2##�2% 3#:B5C#:BES#:B Uc#�"e� 4t�&v��2xk[ 46�A��Q�P<J��D�A\Ւ��HIS}�zk[� �� 20�21-04-21��V��� 9 +�>_P_b_t_�_�_x�_�_�[L[SQ�18-02-27�_�_ok@��; Đ�B�b;c!�DQo�couo�o�o�[ZB���X6�_�o�o#o :���s.@Rd\v�ZY���X5�o����������B  7 ��p� 8 �:�97 �2d��Ko�ZTI��X�"�����l����I��@: ��������(�:�LS���W19��n���H������h�A6`pBdxtF�Ea�:d9�Db㕗S���XPK& Q��oI�[�m�9�9bF`K&Cc������ʯܯ���M� �O_;��7+P[�c�u������� ��Ͽ��_�_?�)�;�$)h��d9`�AdA`Y� I`Y�DχϙϫϽϫo@�o���)hqdp 5� �S�e�w߉ߛ߉ ���������+�=�T+���c9�8'P_A�Y�I�83�^Q�a�D� k�}�������ŏp�� �1�C�U�C�U���� ��������a�ѐY�ِ 5��Y��a�9�Y��� y�2 �2���z�z� Y������������ �&�`%PT ��������//�]J/\/%lBҁ�C7!f�DjC E i/�/�/�/�/�/��9/ &?8?%l1bpAE?t? �?�?�?�?�߼�?O@O(O:OLO^O'��19�#�1f� I�1bQ� 1b�O����O�O�O�� _4_F_X_j_|_ j�|��_�_�_�_�_Ö�Qѐb��b�b  b9�b��bJo\o@J\�o�o�o��a ���b�o�o&8�&I_CFG 2�{: H
C�ycle Tim�e�aBusy>DwIdlzr�t�min={�q�Upvv|qRe�ad�wDow��x�ۂqsC�ount|q	Num qr�s�={��`y�q�PROGWr[|:D�0� u���������Ϗ�y ��SDT_ISOL�C  :�r��?J23_DSP_EN~ �>#�?INC }��e��A   ?�=���<#�
�>j�:�o u���`���a��ȟ�OBK��C,�FeU��G_�GROUP 1~��< A� �j�Cy.�П?Dxd�m��`Q�������̯�����&�Dw���ڙG_IN_A�UTOdQ�#�PO�SRE���KANJI_MASK���t�KARELMO�N :(��by ���(�:�L�@~²JO��V�X��nż����CL_Ld�N�UM0�����EYLOGGING`�?�j�U�F�LAN�GUAGE �:
��DE?FAULT �(�LGXq�V��r��d�  8԰p� ��`'�G  ɤ�`�ۏ�;���
��(UT13:\\Ϧ� �ߵ� ���������!�8�E��W��(��#LN�_DISP ��M��x������OCT3OL���aDz@���f��GBOOK �)ݹz�qz�z�� Xr�k�}������������5Ӱs����	-�t�*��/ُ`��+�_BUFF 2��� A2 �uv�ꂒ�w�� ���#,YP b���������/��ZDCS �V�Y�n���#Dx�^u�/�/�/�/6$IOw 2�B+ cp�/cp@���/??*? >?N?`?r?�?�?�?�? �?�?�?OO&O8OJO�^OnO�O�O�O�%ER/_ITM��dD��O _#_5_G_Y_k_}_�_ �_�_�_�_�_�_oo�1oCoUogo	��BSE�V�����FTYP���O�o�o�ovm���RST��4%SCRN_FL 2��-@��g/gy��0���TP������b�NGNAMp,�`�
�2$UPS��SGIp��U�B��_LOAD�G �% �%DRO�P��MAXUA�LRM�®� �rU�
��H�_PRM���� !���C����7������Pw 2�7� �q�	�ol�W���{���Ɵ ���՟���D�/� h�S�������¯��� ɯۯ��@�+�d�v� Y�������������߿ ��<�N�1�r�]ϖ� yϋ��Ϸ������&� 	�J�5�n�Q�cߤߏ� �߳�������"��F� )�;�|�g������� ���������T�?� x�c����������������DBGDEF ���[!��_L?DXDISA-��{��#MEMO_AP�'�E ? �
 $x(�����������FRQ_CFG ��m(A x'@�E��<[$d%mt$:������*�/� **:�����_ ����+/"/4/a/X/ j/�/����/�@�/�/�/�/�',(�/>?�$ ,?i?P?�?t?�?�?�? �?�?OOOAO(OeO�wO^O�O��ISC 31� �� ����O ��)�O��2__V_�O��B_MSTR ���myUSCD 1�o�N_�_J_�_�_ o�_4oo1ojoUo�o yo�o�o�o�o�o�o 0T?xc�� �������>� )�N�t�_��������� ��ˏ���:�%�^� I���m�������ܟǟ  ��$��H�3�l�W� i�����Ư���կ� ���D�/�h�S���w������Կj_MK'�]Y�$MLT�ARM&�-� 3" P�X�> METPUK ǲ����YNDSP?_ADCOLr�& �}�CMNT�� Ɔ�FN���τ�FS�TLI���ǁP ��^'�G�Y?�IԆ�_POSCF�����PRPM��Y�STv��1��[ 4Q#�
��ϱ������ ��������7��+�m� O�a��������������E�/��SI�NG_CHK  }��$MODA%���K���DE�V 	N
	M�C:��HSIZE�Kǰ��TASK� %N
%$12�3456789 � 2}�TRIG ;1��[ l^�9n�=YP���5��~�EM_�INF 1���`)AT&F�V0E0�+)�E0V1&A3�&B1&D2&S0&C1S0=)ATZ+f�H��:��bA��/�'//K/]/  �/5GYk�/�  ?7/$?6?�Z??~? �?w?�?g/y/�?�/�/ �/2O=?�/hO�?�OGO Q?�O}O�O�O
__�? @_�?OO)O�_MO�_ �O�_�_�Oo�_<oNo 5oro%_7_�o[_m__ �o�_&]oJo �;�����o� �o�o�o�oX�|��� ���e֏�����|0���NITOR��G ?��   	EXEC1˳�s�2y�3y�4y�5�y�C {�7y�8y�9˳t��rޔx�ޔ�� ޔ��ޔ��ޔ��ޔ���ޔ��ޔ̒ޔؒޓ2��2�2��2	�2��2!�2-�29�2�E�2Q�3�3�3����R_GRP_�SV 1�  �(7񿩕�?����0B��r�;T�ǯo@�3S&��
_Dς��~9�ION_DB������Ǳ  ��������~���q�싷�  �ī�Ŧ�&�N  W ������ h�� G��-ud1�����υ�PL_NAME !�<��!Def�ault Per�sonality� (from FsD)����RR2��� 1�L6�L�A�<��� d:҉ϛϭϿ����� ����+�=�O�a�s� �ߗߩ߻����������2��.�@�R�d�v�@��������<� ����0�B�T�f�x�����������޲�D����
���P J\n����� ���"4FX '9������ �//0/B/T/f/x/ �/�/k}�/�/�/? ?,?>?P?b?t?�?�?�?�?�?�?�> �H�6 H�b �H\���  �O1M�dC@PO bMFO�O�G@�=�|C��O�M�O�O C  �H__ _2_P_V_t_@�_�f��_�\��E�	`_�_o o�Q:�oA`�@oRodo�vn A�   �i�O�o�Lޱ�o�k�O �o'9$]H�:J�R�� 1�4ɴ���R@ � �&�<��p @D��  �q?��s�q?���q�A��6E�z  �q���;��	l�r	 ��@� �0�ް!� ���p� � �� �F��J���K ��J˷��J� �J�4�JR�<g|v�f0O����@�S�@��;fA6A���A1UA��X{����=�N���f������T;f��X���ڀ��* � ��  �5'��>��p�H���?��?���{#�����ԏur`�f��q{��g�������i�V����(  ����¤��Ȗt柉�	'�� � �I�� �  ���e��:�È(�ß�=���@���߶� <!��� � �  ��qz�˂�r�o�o����ү � '覵��@!�p@�a�@���@��@��C�C�"��"��B�pCz%����@�r��������n���� ���m;a;n�`@����D�u՟ҿ����῀��Q�c�E�UŔ��w :�W  x�x?�ff�O�Ϙφ*� �P���ˍ�8x�����>��x��q����0�P:�U�7�x0�0���>���|����<2�!<"7��<L��<`N�<D��<��a,h��ߴ��s��s| ҈`?fff?���?&�аT@T����?�`?U��?X�ᒩL� ���t,��t8��wW��� ��ό�w������ �����.��R���!�F��A���=���)����M����HmN� H[���G� F��HZE ~i������ � �oAK���� ����)���/ ��%/7/�j/U/�/y/�/�/��M��"�i���C�/?�/5? =8��`??F??j?��ç�sY��-M�BH"��.��?,�[2�Y0X1�1�@Iܔ=@n��@��@:� @l��?٧�]�? ��%��n�߱����=�=D���0OB@��@��oA�&{C/�� @�UXO�+�J8��
H���>��=3H���_�O F�6��G��E�A�5F�ĮE���O�@��fG���E��+E�?�EX��O�@�>\�G�ZE��M�F�lD�
�p�O�?E_0_i_ T_�_x_�_�_�_�_�_ o�_/ooSo>owobo �o�o�o�o�o�o�o =(:s^�� ������ �9� $�]�H���l������� ۏƏ���#��G�2� W�}�h�����ş��� ԟ���
�C�.�g�R� ��v��������Я	� ��-��Q�<�u�`�r����fB(hA4�̯�h���൘�3��ϩп��!4 ��{����!�0+#8(�:��jbT�f�1E�䴛|�� �ˀ��Ϯ��������JiP��P:�IV c߶�oߙ߄߽ߨف����������9�$��"$<�N��r�����v�H���&��e ,�6�l�Z�|�����n)���������8F
  2 H��6�&H�{�g\Ŵ�&B�!�!� B��0�0A� @�/��$��3����l ^pUgy���$�0� � ��r� T�%
 � �//+/=/O/a/s/ �/�/�/�/�/�/^J�� ��$����4��$MR_CAB�LE 2�$�� � V�TP�
�@n�?�0F1�?0S��0z Bz C[0�n�OM�`B��^��R6>n�:n��F���n�??Q6�  B�� TO�
�vr0��&���n�n�E��O�|Œ?�8� �� C�� 9h4��r0�^��.�~n��2g9y��?�?�*\0��� [@CW@j27�(�1n�=xP�2I�/T3�OR˰O�O �O�O�O_�O�O"__ *_�_�_`_�_�_�_�_(�_or5 +��_Qo couol�?o�o�o�ol�w*�o** 3�OM �%9���zn���%�% 234567O8901%7u "PRFqn�[@ �n��n�
Lw�nn�ot sent ��jzsW,�T�ESTFECSA�LGRI�gkʝd��t��q
�tG �P�n��"��'�9��K� 9UD1:�\mainten�ances.xm�lS���  ���DEFAUL�T2GRP 2=�	z  p�S�n�  �%1s�t mechan�ical che�ckL}n��6��>�G�H�$r����������n��co�ntroller ��7��Ic�8�`J�\�n���ϑM�,��n�"8��n�ȡϯH'�����*�<���Cٟn�����Y����ҿ����ϒ�C�ge�. b?atteryς�W�H	���ϖϨϺ����ϑSupply greasK�,��È�
�<���Hs�H�Z�l�~����ϑ �cabl��߾�g�
7��� 0�B�T��ؑ+�����Q������������`�$��@�hoo�  �����������+�  O�a�s�)Zl~� ����'9  2DV���{ ����
//k@/ R/�v/��/�/�/�/ �/1/?U/g/<?�/`? r?�?�?�?�/�??-? OQ?&O8OJO\OnO�? �O�?�?�OO�O�O_ "_4_�OX_�O�O�_�O �_�_�_�_�_I_om_ _To�_xo�o�o�o�o o�o3oEoWo>P bt��o��o ���(�:���p� �_����ʏ܏� � O�$�6���Z���~��� ����Ɵ��9�K� � o�D�V�h�z���۟�� ����5�
��.�@� R���v�ůׯ����п �����g�<ϋ��� r����ϨϺ�����-� �Q�c�8߇�\�n߀� �ߤ������)�;��� "�4�F�X�j�ߎ��� �����������m� ��T���C�������� ����3�i�>�� bt������ /S(:L^p��	 T~�� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�?�OO0OBOTOfOxO � �?�  @� ��O�O��O��O__(_�;*H_** �� �@zO|_�_�_b_�_�_�_�_��!__ �_Ko]ooo1o�o�o�o oo%o�o#5o Ak}��o�oQ� ��E�1�C�U�� ��a�����ӏ�����	��e�w��
�$M�R_HIST 2���v�� 
 �\�$ 2345?678901����P�BR��9���� �����?�Q�c��,� ������t���ԯ�� ί;��_�q�(���L� ��˿��￦��%�ܿ I� �m��6ϣ�Z�����ϐ���[�SKCF�MAP  ��y��B������ONREL  ��v�.�6���EXCFENB�`�
,��y�FNC���r�JOGOVL�IM`�dv����K�EY`�����_�PAN_������R�UN����SFSPDTYP��k���SIGN`�r�T1�MOT��o��_�CE_GRP 1��.�~���O ��÷���a������ C�U��y�0�����f� ������	��-?& c����t� ���Mq�(�QZ_EDI�T]�(�Q�TCOM_CFG 1�$�a����� 
�__ARC_}�`����T_MN_MO�DE]���UA�P_CPL/��N�OCHECK ?�$� ��  �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�?�I�NO_WAITc_L\���NT���$�3���1_7ERR��2�$�6���OEOWOiO�L<юO��O�53 OC�#M|� C�f���Bvſ��ԹX�²�_C~���<�� ?���_�O?�|7NBPARAMB]�$���Df��_b8ѫ_�[ =  ���_�_�S�_o(oo 4o^opoLo�o�o�kb���o�l}_n#U�M_RSPACE�!��b�GQt�$ODRDSP#_���OFFSET_C�AR�_/�vDISܑ�sS_A3 AR�K]�OPEN_FILE�p_����cqPTION_I�O�����M_PR�G %3z%$*�A�S��sWO�p����C쀄���.�  ;�?֞�9�g��	 ��Ȟ�ڵ��4�dpRG�_DSBL  �n�.�J��sRI_ENTTO_����C�>�-�A �rUT_SIM_D��+ҋBdpVhpLCT ��=���O}z��d\�_PEX; ܳ��RAT;' d�����pUP )�m��pw����� �>�L��$PAL��2��>`�_POS�_CH�p��`�ZP2���L6�L;A�W����o ѯ�����+�=�O� a�s���������Ϳ߿@���'�9ϵ�2�� h�zόϞϰ������� ��
��CW�4�F�X�j� |ߎߠ߲��������� *wS$�4�5�4�Z�
BPG��������� ����&�8�J�\�n� ����a�s��������� "4FXj|� �������� 0BTfx��� ����///_��g�Y/k-���c�� �/�+�/�/�'>->-�o?�/3?�'tP(7R? H?Z?l?�?�?�?�?&0`w��?L�D(4	`<?�6OHOZOA:�o�<�xO�O�O�O�`A�  �I!?�O�__ �]?>_)_b_M___�_��_�_u����O�1������ ��$B@ ��؄��P @D��  a?�c�Q?�<�a<�D�  E�z0c�:�;�	l�&b	 �@�� 0�PP_` �
`�� � � ���b�PH0#H���G�9G��ģG�	{Gkf���GΈK/�o�l�P�C�1��`[�D	� D@ D7g��n�d���  ß5��>(p`�p4�(: B4��Bp{�!�<���O��" ��r'a�sW�Ao�R�ҧpߐ�p(�  ��p�����_$��E	'� �� B�I� ?�  ��E�F�=���f�x��߶� <_`�� � � ��ف��8�" b__�GN=���  'N�(��aOpC��`��`[pB`C�c5�G� ���@��i���~�m����G�MuAuN�@@<��*b 7e����4��X�C����������<�� :��a�tx?��ff�/į֯h� @��O�8<�3�A�>�׶q"a�J�pn�Px���uancnd؃�>������u<2��!<"7�<L���<`N<D?��<��,�o㿌�c� c^��@?offf?�?& ���D@T�2�?��`?Uȩ?X�B�:銒�'d�I ev�g���Zd���� ���������6�!�Z� l�Wߐߢ�y��߱����aσυ���D���Hm�N H[�ArG�� F��M��� �����������(� �%�^� _���K�� ���+���g�*< N�cu������Β���I�={C�O�s^?��}���?yKç'c�'sqH�`E�xp��������:!@I�>}@�n�@��@�: @l��?�٧]/ ���%�n�������=�=D���n/� ��@��oA�&{C/� @�U�/� �+J8���
H��>��=�3H��_�/ �F�6�G���E�A5F�ğ�E���/� ���fG��E���+E��E�X�?� >\�G��ZE�M�F?�lD�
`8? /�?n?�?�?�?�?�? �?O�?OIO4OmOXO �O|O�O�O�O�O�O_ �O3__W_B_{_f_x_ �_�_�_�_�_�_oo -oSo>owobo�o�o�o �o�o�o�o=( aL�p���� ���'��K�6�H� ��l�����ɏ���؏ ��#��G�2�k�V���@z�������韤"(�!�4�ퟦ���<�֕3�ϩ� ��!4 �{:�L��!��0+#f�x�Z��jb����1E����|�������쯠"��F�4���P޲Px�����������׿¿��湿����A� ,�Q�w�bϝ"$zό� �ϰ�����ߴ���@�.�d�R�ej�tߪߘ�0��������)�����.��R�@�v��  �2 H�6�&HY�����\��&B#L#B�  A� @'�����"�4�F�W���߁�������������$�� �� q�� ��%
 ��3EWi{ ���������* ��b�����4�$PAR�AM_MENU �?����  DE�FPULSE�+�	WAITTMO{UT�RCV�� SHELL�_WRK.$CU�R_STYL��OPT���P�TB��C�R_DECSN�i�<, 6/H/Z/�/~/�/�/�/ �/�/�/?? ?2?[?�VSSREL_IOD  �����j5�USE_PROG %e%W?�?k3CCR�|2��m�7�_HOST !Fe!�4O�:T���?-C�?A/CiO�;_TIME�|6�5�VGDEBUG�z0ek3GINP_�FLMSK�O�IT�R�O�GPGA�@ 2�Lp� [CH�O�H�TYPEbn� V?P?�_�_�_�_�_�_ �_oo?o:oLo^o�o �o�o�o�o�o�o�o $6_Zl~� �������7���EWORD ?	�e
 	RS��@�PNS���s�JO!�TyEP@}�COL�h3���3WL�0 ��՜	���5d�ATR�ACECTL 1��o .v�U V������|&���DT Q����S��D � 7t`�	 �f�$Pf� f���f�v� ����	��
�d�u�ᦒc�uj�u�r�uz�u��	���R����c�vj�vr�vz�v��t��a�s� ��������͟ߟ�� �'�9�K�]�o����������|0���������������! ����䡃2 ��,�>�P����� Ưد���� �2�D� V�h�zόϞϰ����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r��0������\� � ������������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�? OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �U���_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����_0�B�T�f�x� �ϜϮ���������� �,�>�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������//�*/</N/X!�$PG�TRACELEN�  W!  �_�V �l&�_UP ������!� �!�� l!_CFG M��%�#V!� ���${#�/�(�-�  ��%�"DEFSPD ��,�U!~ �l IN~� TRL ��-��!8�%C1PE_C�ONFI� ��%O��!�$�)�l LID�#��-	~�9LLB 1�~7 ��$B�  B4�3�& �5JOE��/ << T!?�1KPO1OHOjO �O~O�O�O�O�O_�O��O_L_2_T_�_�Z B�_�_�_�_3O�_"o�o'oXo�9GRP �1��<W!@�  �[�V!A�?x�D P�DV�C2�� o�V d,D�i�i�1�0��0Wo)O�1�n#´(s
�kB+pRq�2.hR�V!>'oY>a�����~� =N�=R��3��0� i�T���x����Տ��x����  Dz0�9�V 
 �a��q��� ������ߟʟ��'� �$�]�H���l������)W!
V7.1�0beta1�$�ܠB(�A�?\)A�G��aޡ�>�������ޡA����f�fޢA�p��AaG��Q�Q@�(��`� ��K�]�o����#Apأ�r�0 ����Ϳ߿ڢU!��} ���v�$��H�2ϝ:�KNOW_M  ��%�&�4SV ���9��5 N�����f�9�$�6�Po��"�m�3Mvc����} ��	�"V ���T���PܽԿ���פ�@1ߠ���(�wPV�1MRvcĥ�T~��D��u����OAD?BANFWD�ϡ3{STva1 1ś)��4�5���� �&��� �Q�D�V�h� �������������� 
O.@�dv������2�����V �<%�w`3 !3E��4bt����5�������6//,/>/��7 [/m//�/��8�/�/X�/�/��MA���d�3�'OVLD � ;�ߊ���P�ARNUM  p��?�?��SCHS9 a5
�7�1�9��
EUPD�?�5uTO>�%_CMP_��V0�����'��lDER�_CHKzE��`��ҎFwO�KRSg����pa_MO���H_��O�%_RES_G
���;
8��oi_\_ �_�_�_�_�_�_�_o �_/o"oSoFo9?+U6\F_xo+Ua�o�o �o-S��o�o�o-S  27-SZ Rqv -S� ���-S 0�x��-RV 1���|���@`z$�BTHR_INRg��X1����dc�MASmSp� Z��MNo����MON_QUEUE ������@����$Nq@U�AN8��ۈ�END��_��EXE ��6@B�E���OPTI�O��[��PROG�RAM %Պ%��.��?�TAS�K_IU4g�OCFG �Տ�?ɟ���DATA����@(�2��k�}��� ����^�ׯ������ʯC�U�g�y�,�IN+FO���I���5� ҿ�����,�>�P� b�tφϘϪϼ����π����(�:ߕ�����I� di���@DIT ���߬���WERFLA�V����RGADJ �^��A�  ��?�@`�w����� ��W�_�?���z�N�@<@�9���%?`h���dm�C�2�%�V��	H�l7�U��2�?G�A ��t$���*��/�� **:���@�����2�5,�'�����1��1W�9�Q����/� A�o�e�w��������� ����]G=O �s����5� �'�K]� ��/����� y/#/5/c/Y/k/�/�/ �/�/�/�/Q?�/?;? 1?C?�?g?y?�?�?�? )O�?�?O	OO�O?O QOOuO�O_�O�O�O �O�Om__)_W_M___ �_�_�_�_�_�_Eo�_ o/o%o7o�o[omo�o�o�oN�	�<��* cNt����Q�M����PREF S�%�����
��?IORITY��܆}���MPDSP������C�U������OoDUCT�������OG��_T�G��钍ڂ�HIB�IT_DOA���TOENT 1Ӊ�� (!AF_�INEm� �+�!�tcp+�S�!�udB�{�!�icmj�qXY��ԉ����)�a ��ߟ����ٟ ���	�F�-�j�Q�c� ����į�������H�B�T�*����%����V����>}5o�f��/	�����һ��~��AG�,  ��o�D�V�Ph�z��պ��Z뿠�������ϻ�i�E�NHANCE )�u�s�A��d�P�7�~����������PORT_NUM�n������_CARTREP�|Ĝ�SKSTAm���SLGS���ě�G�T�Un?othingX�5��G�Y��{��TEMPG ڑ�e��e��_a_seiban���������"� �F�1�j�U���y��� ����������0 @fQ�u��� ����,P; t_������ �//:/%/^/I/[/�//�/q�VERS�IL����  disablej��m�SAVE ����	2670H�755�(�/E?!`@�G?Y?|�}? 	�8Hw��o�;�?��e�? O"O4OFOTJ�<|?�O��5_�� 1�
ě20�@r�e�Ox�O�g�pURGE�1B掘�WFP�p����W�3T�ѯ��WRUP_DEL�AY ���&UR_HOT %!v�z�?߳_DUR_NORMAL�X���_�_�WSEMI�_�_;o��qQSKIP�C�|��Cx�/�o�/�o�o �o�m}�o's�o!3 EiW���w �����/��S� A�c�������s�я�� ����ߏ�O�=�s� ����]�����˟��|�SRBTIF4T���RCVTMOU������/�DC�R�C�^i �ЗaB4��B��q(B[k@���k?�5�* ��{�m����#���A�ߒ���� $����oۯ�o <2��!<"7�<L���<`N<D��<��9��O֯?�Q�@�u��������� Ͽ����)�;�o��RDIO_TYP�E  �M1�G�E�D�T_CFG ���KbBHSE���Xa2�� �ȸ�����.� � үD�/�h�S��ϙ�(o ���o��ӟ�����;� )�_�M��m�ߴ�9� {��������%��5� 7�I���������a� ������!E3i �����a�]�� �A/e�� �mG���/� +//O/qv/�/G/�/ C/�/�/�/�/�/'?? K?m/r?�/S?�?�?�? �?�?�?O�?!OW?}?�nO;���INT 2��Y���_�G;�� �O�K�+��OX�f�0 _[3O6_'O F_H_Z_�_~_�_�_�_ �_�_o�_2oo*oho Vo�ozo�o�o�o�o�o 
�o.@&dR� v���������<�"�`�N���!�E�FPOS1 1�~d�  x\O ҉���O����+�ŏ ׏�r�]���1���U� ޟy�۟���8�ӟ\� ������-�?�y�گů ����"���F��C�|� ���;�Ŀ_������ ���B�-�f�ϊ�%� ��Iϫ����ߣ�,� ��P�b����Iߪߕ� ��i��ߍ����L� ��p���/����e� w�����6���Z��� ~��{���O���s��� �� 2����ze �9�]��� �@�d���5 G���/�*/� N/�K/�//�/C/�/ g/�/?�/�/�/J?5? n?	?�?-?�?Q?�?�? �?O�?4O�?XOjOO OQO�O�O�OqO�O�O _�O_T_�Ox__�_ 7_�_�_m__�_oo >o�_bo�_�o!o�o�o<Uc��2 1崏^o po�o(LRop �/��e��� �6����/���{� ��O�؏s�������2� ͏V��z����9�K� ]���������@�۟ d���a���5���Y�� }������ů��`�K� �����C�̿g�ɿ� ��&���J��n�	�� -�g��ϳ��χ�߫� 4���1�j�ߎ�)߲� M���q߃ߕ���0�� T���x���7���� m�������>����� ��7�������W���{� ��:��^��� �ASe� � $�H�li� =�a��/�� �/h/S/�/'/�/K/ �/o/�/
?�/.?�/R? �/v??#?5?o?�?�? �?�?O�?<O�?9OrO O�O1O�OUO�O�o�d3 1��o�O�O�O U_@_y_O�_8_�_\_ �_�_�_o�_?o�_co �_o"o\o�o�o�o|o �o)�o&_�o� �B�fx�� %��I��m����,� ��Ǐb�돆����3� Ώ���,���x���L� ՟p�������/�ʟS� �w����6�H�Z��� ������=�دa��� ^���2���V�߿z�� ����¿��]�Hρ�� ��@���d����Ϛ�#� ��G���k���*�d� �߰��߄���1��� .�g���&��J��� n�����-��Q��� u����4�����j��� ����;������4 ���T�x� �7�[�� >Pb���!/� E/�i//f/�/:/�/�^/�/�/?�OT4 1�_�/�/?�?m? �?�/�?e?�?�?�?$O �?HO�?lOO�O+O=O OO�O�O�O_�O2_�O V_�OS_�_'_�_K_�_ o_�_�_�_�_�_Ro=o voo�o5o�oYo�o�o �o�o<�o`�o Y���y�� &��#�\������� ?�ȏc�u�����"�� F��j����)���ğ _�蟃����0�˟ݟ �)���u���I�үm� �����,�ǯP��t� ���3�E�W����ݿ ϱ�:�տ^���[ϔ� /ϸ�S���w� ߛϭ� ����Z�E�~�ߢ�=� ��a����ߗ� ��D� ��h���'�a���� ���
���.���+�d� ���#���G���k�}� ����*N��r �1��g���8?045 1� ;?��1���� ��/�/Q/�u/ /�/4/�/X/j/|/�/ ??;?�/_?�/�?? �?�?T?�?x?O�?%O �?�?�?OOjO�O>O �ObO�O�O�O!_�OE_ �Oi__�_(_:_L_�_ �_�_o�_/o�_So�_ Po�o$o�oHo�olo�o �o�o�o�oO:s �2�V���� �9��]��
��V� ����ۏv�����#���  �Y��}����<�ş `�r������
�C�ޟ g����&�����\�� ��	���-�ȯگ�&� ��r���F�Ͽj�󿎿 �)�ĿM��q�ϕ� 0�B�Tώ�����߮� 7���[���Xߑ�,ߵ� P���t��ߘߪ߼��� W�B�{���:���^� ��������A���e�<K]6 1�h� $�^����� �$�� H��E~�=� a�����D/ h�'�K�� �
/�./�R/�� /K/�/�/�/k/�/�/ ?�/?N?�/r??�? 1?�?U?g?y?�?O�? 8O�?\O�?�OO}O�O QO�OuO�O�O"_�O�O �O_|_g_�_;_�___ �_�_�_o�_Bo�_fo o�o%o7oIo�o�o�o �o,�oP�oM� !�E�i��� ��L�7�p����/� ��S�������6� яZ�����S����� ؟s����� ����V� �z����9�¯]�o� ������@�ۯd��� ��#�����Y��}�� ��*�ſ׿�#τ�o� ��C���g��ϋ���&� ��J���n�	ߒ�x���7 1��?�Qߋ� 	���-�3�Q���u�� r��F���j����� �������q�\���0� ��T���x�����7 ��[��,>x ����!�E� B{�:�^� ����A/,/e/ / �/$/�/H/�/�/~/? �/+?�/O?�/�/?H? �?�?�?h?�?�?O�? OKO�?oO
O�O.O�O ROdOvO�O_�O5_�O Y_�O}__z_�_N_�_ r_�_�_o�_�_�_o yodo�o8o�o\o�o�o �o�o?�oc�o� "4F����� )��M��J������ B�ˏf������� I�4�m����,���P� ��럆����3�ΟW� ���P�����կp� ��������S��w�����6����߷�8 1���l�~���6�!� Z�`�~�Ϣ�=ϟ��� s��ϗ� ߻�D����� �=ߞ߉���]��߁� 
���@���d��߈� #��G�Y�k����� *���N���r��o��� C���g��������� ��nY�-�Q �u��4�X �|);u�� ��/�B/�?/x/ /�/7/�/[/�//�/ �/�/>?)?b?�/�?!? �?E?�?�?{?O�?(O �?LO�?�?OEO�O�O �OeO�O�O_�O_H_ �Ol__�_+_�_O_a_ s_�_o�_2o�_Vo�_ zoowo�oKo�ooo�o �o�o�o�ova �5�Y�}�� �<��`�����1� C�}�ޏɏ���&��� J��G������?�ȟ�c��ҿ�MASKW 1���0��>��XNO  ��=�C�MOTE � _�  ��_C�FG 휭���PL_RANG蘡����٦OWE/R ������SM_DRYPRoG %��%���I��TART ��	�W�UME_P�RO&�8����_E�XEC_ENB � ����GSP�D��ΰָ�T3DB��RM���I_AIRPUR�� ��m�p��M�T_�T�����O�BOT_ISOLEC]��l�̥ȥ��NAME ������OB_OR�D_NUM ?�	�i�H755  ��@�R��d��PC_TIMoEOUT� x�oS232��1�`��� LTE�ACH PEND�AN�б�С��������Mai�ntenance_ Cons�������"�ߒ�No Use�����@�R��d�v�����NPO�f���С��ޙ�CH_L���̝��	���!OUD1:1���R��VAIL!ц��������SPACE1� 2�`�
���ХЩ�巓ΦТ��m���< ���?�Y�Y���K lC�|�������� �%<�Qr Y`�d������ Y)/@/�U/v/ ]/�/������/ /7/-?�/Q?r?�?k? �/�/�/�/�/�??3? )OJO	O_O�OgO�O�? �?�?�?�?OOAO7_ _[_|_�_e_�O�O�O �O�O�__=_3oToo u_�oqo�o�_�_�_�_ �oo)o/Moe� ]o�o�o�o�o� %G=�^����{� ��������!�S� 9����o���g�����:��2��� ��ݏ ����%�W�Z���:� ������Ưǟ3ڟ� ���"�ԯF�x�{���@[���ҿ����4�� ��1�C���g����π�|��������	�5 �.�@�R�d�߈Ϻ� ��ߝ������)�*�6=�O�a�s߅�7�� ����$���5��J�K�7^�p����X� ������E���5V-kl�8��������� y�� f VwxN��G ��� �ń
� �  �// 1/C/U/g/y/���-@���/m�/ȁd0 �/2?D?V?h?z?�? �?�/�/�.�:�?�;O ??�?ZOlO~O�O�O �O�?�?�?�?O_5_ (O:O�Oz_�_�_�_�_��_�O�O�O _"_4o; `� @Ȁme@�/{oW__Y�a�UDo �o�o�_�j�o�o1C aI��gq� ������Q�c� ��7�i�����������Տ�ُ�\
�ol���A��*SYST�EM*�V9.1�0185 ��12�/11/2019� A �� ��r��ӓSR_T �  � $ĐE�NB_TYP �  $RUNNER_AXS� �$HAND_L�NGTH�`�T�HICK��FLI�Pґ�`$INTFERENCE�>�IF_CH���I֑$�9�IND�XD�ĐG1POS?   W�N��`�ANG`�x�_�JF��PRM`�� 	�RV_DA�TAƑ  �$��ETIME } ��$VALU�����GRP_ �  ��A � 2 �SC�ő	� �$�ITP_�� o$NUMڠOUِ�	�TOT�
�DS�P!�JOGLIM�� $FINE_oPCNT@�CO���$MAX�T�ASK@�KEPT�_MIR=�]�PR�EMTq�}�APLD���_EX�������t�@��PG��B?RKHOLD�!�:�I_�  ڲ@����P_MADE��w�BSOC�M�OTN�DUMM�Y163�SV_CODE_OPM��SFSPD_OVkRD��R�LDL¶O�ORZ�TPӐL�E[�F!�[�:�OV�=�SF��ᐓ�T�Fx��A�a�UFRA���TOOL@�LCH�DLYW�RECO1VK��:�WSs�:���=�ROM��I�_\�ڐ @��S���NVERT�OF�S;�CǠD�FWD�t���p��ENAB,��7�TR��`����E_FDO��MB�_CM���B-�B�L_Mi�]��Ҫ�2�S�VSTAA�$#UP�����G�׸�AM����а��%� �3_M��A�AM�A��1�T$CA0�,�D:�7�HBK���VL�IO?�[�IQ�$PPAO�{�`����s��s�1�DVC_DB��F��������A���1��%���y3��+�ATIO� �h�K�U��/�/�P�ABF�T֒E�G��Ԛ���E�:�_AU�X�SUBCPU<�G�SIN_7Ў����P�1������FL�A��ݑHW_C1����j�����$A�TR���$UNI�T�����ATT�RI���G�CYC=LC�NECA!��FLTR_2_F�IR�TARTUP�_CN`Ӷ�SIG�NO�LPS�2�1�_�SCTz�F_��F1_��t��FSF����CHA��[���O��RSD/���/��P��s�_T��PRqO�|�p�EMP�D=��T���ܐ����'DIAG�R�AILAC��p�MF�LO��'�4�PS-�@� i�+�%��PR��SB�  ��C�� 	^$�FUNC���?RINS_TB���=�o�RA��`��7��a�E��WA�Rq�8�BLCUR��$A+	((D�A��G(#%LD@=�?�h�o#��t�o#TI��%�ܐ�$CE_RIA_[SWA�AF��P^���#��%T2\C9K��CMOI��֟DF_LE�_�PmD�"LM��FAПHRDYO��E�RGt H� z���O 5MULSE� ���\0��$JW�Jr���ǂ�FAN_AL�MLV�Î1WRN�5HARDאO�_�O,� �2�1ST�O�Ƶ_���AU���R�(���_SBR���5.�J����CMPINFڐp��-De!8CREG@��NV0l�$�۱DA7L_N��FL����$M 2��7%�ܐY�8�ECM-�N0��Y����G���vSP$R�$Y���Z�� �ۡ��7� ���EG!`
��?�
QAR�0�'�2p0�U3 ��AXE$�wROB!�RED!��WR�߱_i]�S�YܰDQᰋVS�WW�RI�V��STRP �)��f�E��Ġ&To�1�B�P1��V�5c�OTOHAĠ�ARY�b]��ΡR�FI��h�$LINK�!��3a?$EXT_�S1��%U6�[aXYZt�2ej7sfOFF9�R2bZbNh`B����d�����cF�I �g�A�7Ĩ9�_JL�¢d�?ch�h�0�T�[8�US�БB	qL2ArC7 ��D�UO�$V9pTURB�0X�#zu!a(BX�P,�)wFL[`��@�P��p|e�Y30�G� W1ĠKF�M�'�3��s�����a�ORQ.���x�� s��m�� �H��,��_A]�OVEd���M h l��C~��C~��B}� �0{�B�|���{�~�� h� ��e�u�����l� v�e�����C���.�SERK��	tE�H���E�A�ܐ�e�� gN!K�N!AX �¢N!���4b��0 ��Z1��o��`��r`����`��:p��qp��1 �p��:0��:0��:0Ǚ :0י:0�:0��:0��:0�:0'�D�8�DEBU��$��3(�N�VbABNL�t�r^�VA�� 
� ���+���7�0�7�o 7�a7�ra7��a7�:q�7�qq�$Fp�"ۂ�cL�AB�b)�����G�RO: )r�<*�B_,��Tm��`�0���*���1�AND �pt�:�+�_e=��1Y� *��A�Pm�!|�- �^`NT�0ӟ�VE�Lل��L���S�ERVE���@ i$�`�A]!���PO@ҹ ��`����¿!�@  �$�TRQ�r
� �tR
���"2��q I_ 	 ql���[ERR�b�oI,��لr�TO	QلրLHP���R��J G��%Ha�� �@��REP  
 �,��#�=�݁RA~�� 2	 d��ps��@��� �@�$r�� ����� �OC?!� � d�COUNT��Q��FZN_CFG	� 4��aF3T������ܣq ��ӼQ��C �(�M ��g2��Ճ{����CFA� 䅻&��XdP@�����SQ��G�rdQPB�"�HEL}@~Y� 5p�B_BAS��RS)R`F�^SS��!RM�1��M�2p�3p�U4p�5p�6p�7p�98��@�ROO�p���V ]`NL�ALsAB���FN�ACK�I%N�Tg �CU�0E0� 	_PUdq�2ZOU��P�aH-���� �P��TPFWD�_KARw�iAf�R�E��$0P/`U!w�QUE`I e�Up�r�0�1I�0�-�[`S��SF[aSEM3��A��0A��STYSO� 	�DI�}㸻���!_TMuCM�ANRQL[`EN�D�t$KEYSWITCH^s.��HEUpBEATmM�PEPLEv�(����UrF�s�S3DO_HOM�� O�1 EFA�PAR�a�vQ�P�EC��O01c���OV_Mxr� � IOCMGt��A����,�HK�A DXabG��	U^ҹMP�W�Ws�FORCfCWAR� 2��.�OMP G @��c�0U�SEP3P1�&�@�$3�&Q4����O� L�"y��aHUNLO9 �\�4ED�1  ��SNPX_A�SZ� 0�@AD�D��$SIZ�fA$VA���M_ULTIP��.3�� A�! � �$H	/0��`BRS�}�ϱCrТ6FRI	Fu��S� �)��0{NFOODBU�P�~��5�3�9�ƽAfI�A�!$V�y�x�R�S|N��@ � L0Ə�TE�s8�:sSG%LZATAb�p&o�sCx᳍P[@STMT�q2�CPP�VBWe�\D�SHOW�Ev�BAN�@TP�`�wqs8���s8��r��V7�_Gv�� :p$PCD X�7���FB�!PX�SP� A U�AD�P��� �W�A00^�ZR� bW@� bW� bW� bW5`YU6`Y7`Y8`Y9`YA`YB`Y� bW��cV�@bWF`X7�$hlY(@�$h�Y@@$h�Y1�Y1��Y1�Y1�Y1�Y1��Y1�Y1i1i1�"i2_Y2lY2yY2��Y2�Y2�Y2�Y2��Y2�Y2�Y2�Y2��Y2�Y2i2i2B"i3_Y�p�xyY3�YU3�Y3�Y3�Y3�YU3�Y3�Y3�Y3�YU3�Y3i3i3"iU4_Y4lY4yY4�YU4�Y4�Y4�Y4�YU4�Y4�Y4�Y4�YU4�Y4i4i4"iU5_Y5lY5yY5�YU5�Y5�Y5�Y5�YU5�Y5�Y5�Y5�YU5�Y5i5i5"iU6_Y6lY6yY6�YU6�Y6�Y6�Y6�YU6�Y6�Y6�Y6�YU6�Y6i6i6"iU7_Y7lY7yY7�YU7�Y7�Y7�Y7�YU7�Y7�Y7�Y7�YU7�Y7i7i7"d���VP�U�# �߰e�
�A�2��� x #�R��@  ��M��RX9� ��Q_+�R��P��(�~ ��S/�C�D�^�_U�0i����YSL���� � L5Bj��4A7��D����&RVALU�j�% x1���F��IgD_L�3��HI���I�"$FILE_L!�i$�� ��{SA� h	�~M�E_BLCK��Z�uAc�D_CPU�s�M0s�A0u�$�6�E����GR  � PW-����06��LA�AS��������RUN_FLG���� ���v�!���!���HF ��C���vl1T2x_LI�"�  ��G_�O�� P_ED�I�"D@T2��c��k�9��nє0�0 ��TBC2LT �Q@ �(0�!c��FT���	TDC"�A4z���M����L���TH�0�!��#�$�R��0e ER�VE�F�	F�5A��� �  Xw -$q�LEN�0~�	q�) RA� 2&��W_?���1q��M2��MOk�5S�0 I. Z�����q����DE�1LACE,":�CC3Z¶_MA20>>GTCVEfTX g
�|
8R1Q�*1QJA-UM��БJ>JP�}�2��@0P	0JKVK�A.)A�.5A#J�AF2J�J:JJBAAL�2h:hbAAf5#� N1��XB 
G�L��_�A�0ٱm�CF62! `	�G�ROU��vA�2$QN���C�3�REQUsIR1��0EBU�3�m��$T 2 �*!n�&��50��" y\� ��APPR  [CLG�
$t�Ng('CLO��w)S��)r
��u6# ����M �C � 2�$_M	GA� CLPN��(� �R �'BRK�)NO�LD�&�@RTMO�b�:
=�%Jb�4P j  :  B  �  �  6W57W5hAn |���$� "Ę��A�7)A�3PATH�7�1�3�1���3� / #\�PSCA��� 7h"�!INp�U�C����0@C:PUM9HY���� @A���L�[J�0[Jq0[@PA�YLOA7J2L��R_AN��CL��ЦI�A�I�A�%R_?F2LSHR@��ALO�D~A�G=C�G=CACRL_��-E P�)G�D�H��G�$yH�"NRFLEXj#u��J��% PT"�����E�W��Z�BJ>p�& :}���  �W�T��� ������F1�QEeYg���� ��(�bE2D Vhz����`x }t��m`�x��H�QT�w^qXF� ��d�h%.�x1 CUgktb��������BJ�' �����	/���cATrf!� EL�`�(�D�#(J/ &* J�E0CTR)AmaT�N��@�'HAND_VBG�jQ���47( $�pF2�&�-��SW��"�&)� $$M�@ �)!��!�1�#p��E2�A���@�&��<���-A�,���*A;A�;G��+���*D;D�;P�0G��ݩST��'�9�N8DY �e �&(�O��@r��G �Q�G�A�G�t`�5P_5h5q5z5�5�5�5�2�J��* ��T�2 �a㵙!��ASYMEZ�� F)K� L�A$O_ B�X5@HD2=4ĸ�ROdOvO�O�CJ�LR0�Jp�����Id_VI���ؙ#!�V_UN ���6�W��AJN� |�N��LR�U_ԃ�]�� $YR03_E_���0[TcS�"��HR����+���}P]"DI�0#O#�2��S, g�V�I9�AV1 SP�s`^�^�v`���`�� - � ɑME�a��y���`�T�PT��Հ�0����V ��������T��� $�DUMMY1q1o$PS_p`RF2`�  �0���PFL�A�YP���?$GLB_T��1���]! ��aq�}��. XT '�1ST��* SBR�0M�21_V�T$S/V_ER�@O��w��CLK�w�A�`OlS� �GL�EW��/ 4���$Y
��Z��W���Aœ�Az�9B肼�U��0� �pN���$�GI��}$�� �/������1� L���}$Fz��ENEAR�`�NwcFd	�`TANyCwb��JOG&`�H0 2�$JOINT�"�� ���MSET�3  "EJ�a�S����1��4� �n`U�a?�* LOCK_FO�@Б�oBGLVt�GLTEST_XMj N�EMP� �r2I�� $U�P��9`#20* ��X1#̐4� X/y�CE�&�y $KAR$qM>%�TPDRA����VEC`�� I�UX2]HE T�OOL9c�V8dR�E�IS3�U�6�z1m`ACH� / 3��O@����3g��% SIZ"  @�$RAIL_BO�XE���ROB�O)?���HOW�WARVQH!��!ROLM�n%ԁ$"p�6 a`�0O_F��!��HTML5��)AͲ��!�15���R�O�R6��"1`�� �ӽ�O�U�7 d��T/�`�J�$�� $PIP*N�p�6"!`�X� �PCORDEaD� 
@� a XT*0�) � �O`� �8 D 0�OB |�N�� �7v1��/�v2܊�P�SYSv1ADqRO� ��TCH�� 9 ,�pENT	�QA_�4�݁@��.VWVA~|�: � �����PREV_R�T��$EDIT�(FVSHWR�Pc�G@�b���D���O�^DW�$HECAD����x@��0C�KE����CPSP]D�FJMP�0L�2P�R�`;�;~0{Q��6I3SO�C��N�E�P���TICK�9c��M�Qu�CH=NY�< @�0�AᅗA_GP&V-&�PgSTY�2!LOK����C"R�P= tk 
#@G�5%$A�=c�SE�!$@D�9`���M��P&�&VSQU�,e�яTERC�ਁP�S�>  o�� �p��q�``O����F{`IZ����PR\0�Db�A0P9U;�Te_DOi�0�XS� K�AXI4s`�#]UR��c@P�O P�6���_��2ET�bP�0	ŐՐ� 
�sPA�����9'[) ��S=R��?l�P� !���/u�Ay�/u*� /s8�/sH�uuj�uuz� uu���u�}���u�|���yC
��}C�}�ϕϸ�Ϲ�-SSC3� o@ h��DS4P̗��SPJࡅAT�x� �UaP�B��A_DDRES�B3@�SHIF�O_2+CHO��1IR����TUR�I�� }A�"CUSTO�d*�V�I>�B�2���8c�
2
ՒV81da~�C \a�8A�rPC�a�P��C���b�bR�6���T�XSCREEx2Dz��QTINA���# Ӕ\P� Q_��ٰE T�A��8b �1��n� ��a�2�b�/@RROS�~ �0�@���dͱUE�DF ����1
�S��1RSMPwgUe0�P����S_��=Ú���ȧ=õaC����o 2E��UEմ�GD���D`GMTJ��Lp��a~�O��
�BBL_ W���~�H ���J�O��V�LE�a�N ��`�RIGHj�B�RD��ہCKGR�����Tf0����WIDTH#T@�b)!��)�UI� E	Y��}�I
2� m VRz6 @aBACKTQh�Ũ���FOS1n�LAB_q?(��yI �$URT!�E���ް��H@� 'J 8��~ _wA�h�R���s(��@U�O�~�KP$����Uv���Ry!�LUM�ØfՀERIV!1R�Ph �L���`GEI�O�`l2&�@LP��bE�Pf�)%�v�3؆�3�  2�U50�60�70�8Ҁ�R��?`h ���� !��S�PKݱUS=R��M <a���1U(�FO�PRI�am  ����TRIP2!m��UNDO;�N `�P �ye`!xe �O�`�P Oc���CaG PT� T��&^�OS��s�R�`F�J��Z�P��������6TACJ�U�Z�Q����ã�5UJ�OF�F([�R_���O)� 1P���;�-Q��GU�1P:��"pV�Q�`��SUB6R����SRT��tS0R}� #cOR ��'RAU(p��T���7r��_&@�DT |1p��8OWNM��4$GSRCQ�Ҡ�PD(<&rMPFIMTl��`ESPPab�� ��eA�������A@
�7U `��WO[p�4�a�PCOP��	$�`O�_- b�1�WA3@CF�� �Z���@l"+� �V�SHADO�W�`��_UNS�CA��ʴDGyD!�1EGAC�8��VCWp`
�W� ,"w1�S$NER�c�Q�#+�C0cDRI5V6f�a_V/P���@m D��MY_UBY��kyV��UR���P�eA�� "P�_MT"LZkBMv]�$�@DEY�3cEX7�^��MU�@1X]�V$��US���`�_R��R��
�R���QG�pPACIN�A�PRG�$�"�`�"��"ң�RE}遚�:�H�"@XS �� G�P��H� �IR��@Y���?�ӱ��	�qaRmEb#SW� _A�!�<�W#B`O��ہA(�^3/rE��UeP�Z;�6HKjRZ���v:�P&q[0%��3EAP�7� j�^5۰I�MRCV
�[ ���OvPMj�C��	p�2��#�2REF6� F�6�1M0���c50�� �:FAJFAKhE�6�?A_ �:�H�;�pS�ЀN'�aa��I�\ �GR�ӵ`�м�POU4W�"VkO W 5U�2��a$Ԑ��C`,�Y���U�2Q{�ՀULj��Z_ CO~��[H EPNTZ�T��U ���V�ђSQPL��U�#�U���W���V�IA_���] �殐HD����$J�O��6��$ZO_UPL�W�Z|p�W!e�QPSp�0�_L=I��$EPEQ��k�a�QǑ΁��΀K��P]m�^� 0贃�a� ��CACHLO:A�d�aI оi��� 1CI`MI�FHa�eT�p�f�K�$HOj��`C'OMM���Ot�w�WӲ�S&�T7 V�P�"@�mr_SIZwtZ� rx!asw�v��MP�zFAI!`5G�4�`AD�y��MRET�r|wGP���> & �ASYN�BUF�VRTD��%�|q��OL�Di_��A�W��PC���TU7#�`Q{0	�EwCCU�(VEM� x�e���gVIRC�q�9�!���%�_DEL�A�#&Q���AG:5�RK!XYZ̠��K!W1��8A��򱦀TN8"IM߁8���|���eGRABB��Yb"�e�_� ��LAS��<��a_GE�e`u�&��;���T/S&N` ���%aI���"ņ�BGf�V5��PK� ǆ�a�WGI��N#�`2 ����`�qq�a+�a�S�p�fN:�0LEX��b�����;��Nq��I? �-|�� |�.$�3����- �"c��b�t�Ŀ��.a�ORD�����иw�RN�d $MPTIT� �C��F��VSF����e a -�[�QK UR61SM!�f+����ADJ�N%�PZD�>�g DƨBaAL�+`�p�AbPERI|s`��MSG_Q9�s$}q�u  ���b��h+�"�g�J`�^3p�XVR#�in��b�T_OVRi��_�ZABC��j�"(;�s/@
�Z]�#�k+�=$L�-B�1ZMPCF��l�H���A����LN�Kc�
����m� $,q�0��CWMCM� C�C����p4P_A+A$J����Dbq�� �� �� ����
D��F�UX���UXE ]!f��	�]��]�o�p��oё���FTFsQ�Ӿ�r1�Zb��n {�}� d�a��YJ`D�� �oY�R�pU�$�HEIGH�#"�?(MP�.A�P���D�p � EX�$�BQPx �SHIYF�s��RVI`F��/B|�0�C`�dT�F {"�������WuD���TRACE��V���K��SPHER>� q ,MP�<)�;��$R�!p�~� ���F�? S�6��S�F��  �S�x�2p������ s���r�����	���U�C�ADC���l6�R   d�� ZD �Qx0C���l�l0�| ʆ6�V��@ 2�F���� D� P�����	�	F� ,:$ZH~l� ������ // D/2/h/V/x/�/�/�/ �/�/�/
?�/??.? d?R?�?v?�?�?�?�? �?O�?*OONO<OrO `O�O�O�O�O�O�O�O __8_&_H_n_\_�_ �_�_�_�_�_�_�_�_ 4o"oXoFo|ojo�o�o�o�o�o�oF��$S�AF_DO_PULSC�G��k�$qp����|k���5qR� �`�XP�+S�S�
������s��tq  ���������*�<�N�`�r�����]�  ��2��Dtqtqd�������rs�� @�������*�܉�� � 6���_ @J�T�Y J���������T D������� �)�;�M�_�q����� ����˯ݯ��~�����M�_�8$��sR�;��f����p���
�?t��Di��q>��  � ���� R�q|ulq���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e�@w�����S��G� ������0�B�T�f� x������������ ��"4FK��b0E�ҳD�ܽ��� ���'9K ]o������ ��/#/5/G/Y/k/ }/�/�/�/�/�/�/�/ ??1?C?U?g?��? �?�?�?�?�?�?	OO -O��QOcOuO�O�O�O �O�O�OLz��!_ 3_E_W_i_{_�_�_�_ �_�_�_�Yoo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������ø��Ǔ�6�H�Z� l�~�������Ə؏ꏀ��� �2�D�V�d�p#�m�����������i�	123�45678ݲh!B!ܺT
z1!���
��.� @�R�d�v�������"� ïկ�����/�A� S�e�w���������ѿ ������)�;�M�_� qσϕϧϹ������� ��%�7����m�� �ߣߵ���������� !�3�E�W�i�{��L� ������������/� A�S�e�w��������� ������+=O as������ �'9��]o �������� /#/5/G/Y/k/}/�/ N�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�/	OO-O?O QOcOuO�O�O�O�O�O��O�O__)_;_BS��]_o_�?�_�_�_�ԚCz  Bp��z   ��2��� } �X
~g�  	��R�2U_<oNo`oro�l��\�+o�o�o�o�o "4FXj|� �������� �oB�T�f�x������� ��ҏ�����,�>��P�b�t����������Qa�R<Ք �˕a  ��������#a#at�  �P#�;���`��$SCR_GR�P 1*P�3� � ���R �U	 ����������Qԑ�U�������ٯǯ ��]ٰ`��C�,�����m��C����lL�R Mate 2�00iD 567�890!`LRM�|� 	LR2D� ���
123	4��Ц�d��hbճ���}�ݣ}��cDԑ����ѡ�	j�4�F�X�j�|τ����H���Ē� }���į������̦<��1��A���e��WV���Vh`,R���  ��B��PƐ�߮��Ԫ�A�P�� c @�0�ժ�@���F�� ?4���H�P�'��ڪ�F@ F�`Q�Y�P�}�h�� ������������ʩ �����J�5�G�Y�k�B�y���������� ��=(aL� p��o�
'������W`�.4�@�4�>�}�4̧@h��n�PȄ�� ��ݣT_��A��H�����aĲ��1 
/1/C/Q*!�f(r/�/S/�P�#
 b�/�/�/� ?�/$?|,4]�ECLVL�Ў�1����>1L�_DEFAULT�F4������0Z3HOTST�Rf=�z2MIPO/WERFE0�Ur5��4WFDOg6� r5=2RVENT� 1M1M1�3 �L!DUM_E�IP,?H�j!?AF_INEf0+O�3D!FTOZN�!O~O!�ϣO ��mO�O!RPC_OMAIN�O�H��O�_�CVIS�O�I��_b_!TPUPP�UY_IdQ_�_!
�PMON_PROXY�_Fe�_�_uR��_Mf�_Fo!R?DM_SRVGoI9g5o�o!R���o�Hh�o�o!
�@M�oLi�o*!R�LSYNC+Qy�8v!ROS� O�|�4e�!
�CEwPMTCOMd�Fk��!	�rOCONS�Gl��Z�!�rWASR�CaoFmI���!N�rUSB��Hn�� �O�Uc���?�d��+���O���s�П87R�VICE_KL �?%�; (%SVCPRG1ןD�	�2�$��3G�DL��4o�t��5��D���6��į�7� ����/�*�97�<���od������ 9����a�ܿ���� ���,��ٯT��� |��)����Q���6� z���6����6�ʿD� 6��l�6�ϔ�6�B� ��6�j���6����6� ��4�6���\�^�
�ܟ ���������.��� ���8�#�\�G���k� ��������������" F1X|g�� ����	B -fQ�u��� ��/�,//P/;/ t/�/q/�/�/�/�/�/ �/??(?L?7?p?�_DEV �9�UT1:|?~�0GRP 2
�5��0�bx 	_� 
 ,�0x? �?�2�?OO@O'O9O vO]O�O�O�O�O�O�O �O_*__N_5_r_�_ �?�___�_�_�_o�_ &o8oo\oCo�ogoyo �o�o�o�o�o�o4 �_)j!�u�� ������B�)� f�x�_����������� ��M�,��P�7�t� [�m�����Ο���� �(��L�^�E���i� �����ܯ�� ���� 6��Z�l�S���w��� �����ѿ���2�D� +�hϿ�]Ϟ�U��ϩ� ��������@�R�9� v�]ߚ߬ߓ��߷��� ����*��N�`�G�� k����������� &�8��\�C�����y� ��������C���4 F-jQ���� ����B) fx_������ ��/,//P/7/t/ �/m/�/�/�/�/�/?��/(??!?^?e3d �e6	L?�?�?�?�?0�?�?OK%�O5O<C���NA�1NE ^OlGVO�OzO�O�O�O �I"O_JI�O4_"_X_ F_h_j_|_�_�O�__ �_o�_0ooToBodo �_�_�o�_�o�o�o �o,P�ow�o@ �<�����(� jO�����p����� ��܏ʏ �B�'�f��� Z�H�~�l�������؟ ���>�ȟ2� �V�D� z�h�����ůׯ���� ����.��R�@�v��� ��ܯf�п������ *��Nϐ�uϴ�>Ϩ� ���Ϻ�������&�h� Mߌ�߀�nߤߒ��� ����.�T�%�d���X� F�|�j�������� *�����.�T�B�x� f�������������� *P>t��� ��d���� &L�s�<�� ����/T9/K/ /$/�l/�/�/�/�/ �/,/?P/�/D?2?T? V?h?�?�?�??�?(? �?O
O@O.OPOROdO �O�?�O O�O�O�O_ _<_*_L_�O�O�_�O r_�_�_�_�_oo8o z__o�_(o�o$o�o�o �o�o�oRo7vo  jX�|���� *�N�B�0�f�T� ��x�������&��� ��>�,�b�P���ȏ ����v���r����� :�(�^�����ğN��� ��ȯʯܯ� �6�x� ]���&���~�����Ŀ ƿؿ�P�5�t���h� Vό�zϰϞ����<� �L���@�.�d�R߈� v߬�����ߜ��� �<�*�`�N���߫� ��t���������8� &�\������L����� ��������4v�[ ��$�|���� �<!3��T �x����8 �,//</>/P/�/t/ �/��//�/?�/(? ?8?:?L?�?�/�?�/ r?�?�? O�?$OO4O �?�?�O�?ZO�O�O�O �O�O�O _bOG_�O_ z__�_�_�_�_�_�_ :_o^_�_Ro@ovodo �o�o�o�oo�o6o�o *N<r`�� �o����&�� J�8�n������^��� Z�ȏ���"��F��� m���6���������ğ ����`�E����x� f�������������8� �\��P�>�t�b��� ������$���4�ο(� �L�:�p�^ϔ�ֿ�� �����π���$��H� 6�l߮ϓ���\��ߴ� ������ ��D��k� ��4���������� ���^�C����v�d� ����������$�	 ������<r`�� ���� �$ &8n\���� ���/� /"/4/ j/��/�Z/�/�/�/ �/?�/?r/�/i?�/ B?�?�?�?�?�?�?O J?/On?�?bO�?rO�O �O�O�O�O"O_FO�O :_(_^_L_n_�_�_�_ �O�__�_o o6o$o ZoHojo�o�_�o�_�o �o�o�o2 V�o }�FhB��� 
��.�pU����� v��������Џ�H� -�l���`�N���r��� ����ޟ ��D�Ο8� &�\�J���n����� ݯ������4�"�X� F�|������l�ֿh� ����0��Tϖ�{� ��DϮϜ�������� ��,�n�Sߒ�߆�t� �ߘ��߼����F�+� j���^�L��p��� �����������$� Z�H�~�l�������� ������ VD z�����j��� �
R�y� B������/ Z�Q/�*/�/r/�/ �/�/�/�/2/?V/�/ J?�/Z?�?n?�?�?�? 
?�?.?�?"OOFO4O VO|OjO�O�?�OO�O �O�O__B_0_R_x_ �O�_�Oh_�_�_�_�_ oo>o�_eowo.oPo *o�o�o�o�o�oXo =|op^��� ���0�T�H� 6�l�Z�|�~���Ə� �,��� ��D�2�h� V�x�Ώ�ş����� ��
�@�.�d����� ʟT���P�ί���� �<�~�c���,����� ����ʿ�޿�V�;� z��n�\ϒπ϶Ϥ� ����.��R���F�4� j�Xߎ�|߲������� ���ߞ��B�0�f�T� ���߱���z������� ���>�,�b������ R������������� :|�a��*��� ����Bh9x lZ�~��� �>�2/�B/h/ V/�/z/�/��//�/ 
?�/.??>?d?R?�? �/�?�/x?�?�?O�? *OO:O`O�?�O�?PO �O�O�O�O_�O&_hO M____8__�_�_�_��_�_�_@_%od_nQ��$SERV_MA_IL  nUd`��JhOUTPUT�YhoP@�NdRV 2�V  g` (�Q4o�o�NdSAVEzlhiTOP10 2�i d j_ 2 DVhz���� ���
��.�@�R� d�v���������Џ� ���*�<�N�`�r� ��������̟ޟ�����U�eYP�oKcF�ZN_CFG �Ugc�d�a��eT�GRP 2�^��a ,B  � A��nQD;� �B���  B4~�cRB21�foHELLW��U��f�`�ou���%RSR��)�b� M���q�����ο��˿ ��(��L�7�pρ�����  ��a%�����Ϗ͓����oP��������Ǫ�2oPd����ɦ�HK 1׫ ߈߃ߕߧ����� ������%�7�`�[�m�������ìOMM ׯ�Ȣ�FTOV_ENB�Yd�a�iHOW_R�EG_UI7�LbIMIOFWDL�����l�WAIT�4���v���t`X�ܡd��TIMX������VAX`��l�_�UNIT3��iL]CQ�TRYX��e�N`MON_AL�IAS ?e��`heo���� �
t��#�G Yk}�:��� ���/1/C/U/g/ /�/�/�/�/l/�/�/ 	??-?�/Q?c?u?�? �?D?�?�?�?�?O�? )O;OMO_OqOO�O�O �O�OvO�O__%_7_ �O[_m__�_�_N_�_ �_�_�_o�_3oEoWo ioozo�o�o�o�o�o �o/A�oew ���X���� ��=�O�a�s���� ����͏ߏ����'� 9�K���o��������� b�۟������"�G� Y�k�}�(�����ůׯ 鯔���1�C�U� � y���������l���� 	��ƿ?�Q�c�uχ� 2ϫϽ������Ϟ�� )�;�M�_�
߃ߕߧ� ��d�������%��� I�[�m���<���� �������!�3�E�W� i����������n��� ��/��Sew�����$SMO�N_DEFPRO�G &����� &�*SYSTEM*ܢ� 	�RECALL ?}�	� ( �}x�yzrate 6�1=>192.1�68.1.15:�6300 .9416 6�l~�;}
!11 ,> P��/� �� �g/y/�/�0/B/T/ �/�/	?/�/�/�/c? u?�?�/,?>?P?�?�? O?*?�?�?_OqO�O �?�?:OLO�O�O_�I�.copy md�:drop.tp� virt:\temp\+O�O__q_ �_O(O�OL_�_�_o �O�O�_�_[omoo�_ �_6oHoZo�o�oo"o �o�o�oi{�o2 DV����� �e�w����.�@�R� ���������Џa� s�������<�N�ߟ� ��(���̟]�o��� ����8�J�ۯ���� $���ȯگk�}����� 4�F�X������ ��� Ŀֿg�yϋϞ�0�B� T�����	�Ϯ����� c�u߇ߚ�,�>�P��� ����*߼���_�q� ��ߨ�:�L������ �&����[�m����6�H�Z������7�!Rfrs:ord�erfil.da�t0Umpback�;_����j|_!Tb:*.*6��P���2x!:\�+�0 �ew�3!a);�� U��
//�� d/v/�/�6/�Q/�/ �/?�/�O`?r? �?��:?��?�?O /'/�/K/\OnO�O�/��/@O�/�O�O�O[��$SNPX_AS�G 2����,Q� P� 0 '%R[1]@��_WY?�C%W_�_f_�_ �_�_�_�_�_o�_7o o,omoPowo�o�o�o �o�o�o�o3W :L�p���� ��� �'�S�6�w� Z�l��������Ə� ���=� �G�s�V��� z���͟��ן��'� 
��]�@�g���v��� �����Я��#��G� *�<�}�`�������׿ ��̿���C�&�g� J�\ϝπϧ��϶��� ����-��7�c�F߇� j�|߽ߠ�������� ���M�0�W��f�� ������������7� �,�m�P�w������� ��������3W :L�p���� �� 'S6w Zl�����/ ��=/ /G/s/V/�/ z/�/�/�/�/?�/'? 
??]?@?g?�?v?�? �?�?�?�?�?#ODT�PARAM �,U6Q �	U�'JP'D�@'H�~D�-PPOF�T_KB_CFG�  fC2USOP�IN_SIM  ,[sF�O�O�Ov@�=@RVNORDY?_DO  }E�E�RQSTP_DSB�NsBU_aX=@�SR �I w� &�@ESTa_�^�T�CTOP_?ON_ERR_;B~�QPTN �E��P�C�RRING_PRM�_�0RVCNT_GP� 2�E�A�@x 	Q_Poh@>owobo�olWVD%`RP 1LI�@�axI�g �o�o�oEBT fx������ ���,�>�P�b�t� ������яΏ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�]�Z�l�~������� Ưد���#� �2�D� V�h�z�������¿� ���
��.�@�R�d� vψϯϬϾ������� ��*�<�N�u�r߄� �ߨߺ��������� ;�8�J�\�n���� ����������"�4� F�X�j�|��������� ������0BT f������� �,SPbt�����bPRG_�COUN�P�D��R�ENBo�M���D/_UPD �1{[T  
 �gBR/d/v/�/�/�/ �/�/�/�/?/?*?<? N?w?r?�?�?�?�?�? �?OOO&OOOJO\O nO�O�O�O�O�O�O�O �O'_"_4_F_o_j_|_ �_�_�_�_�_�_�_o oGoBoTofo�o�o�o �o�o�o�o�o, >gbt���� �����?�:�L� ^���������Ϗʏ܏ ���$�6�_�Z�l� ~�������Ɵ������_INFO 1=@%& H�	 �c�N���r��@
U�@CIy�=��t����Bvſ���X�n²��C~�⒭>��� @g� A���`=�` >�`� >����� C	���	�(>B��hC3���9!C2������@�D�"(>�N���a�3�]���2���YSDE�BUG�A ��d�))Q�SP_PAS�S�B?c�LO�G =�J! � ����  ��%!�UD1�:\��#���_MPAC��@%�#�@!̱�A� @!�SAV ���y���вC��׸SV�TE�M_TIME 1���K  0 7 $��$C�%��C�+��MEM�BK  @%%!ะ��%�7�G�X�|& � @G����iߎߞ�b�����,��^� y�@��� �*�<�v�T�f�x������� ������� 
��.�@�R�d�v��e������������ (:L^p�������� ��SK�����@RdZX�� "�2s���`�� ����� ����%/7/I/[/O�u$� �u/��ߴ/�/0�/���/��?'? 9?K?]?o?��s?�?���?�4^�?�?�?OO /OAOSOeOwO�O�O�O��O�O�O�O__)�T�1SVGUNSP]Dy� 'c��4P�2MODE_LI�M ��g�0T2�=P]Q��/UAS�K_OPTION�X��g��Q_DI.r�ENB��c��Q�BC2_GRP 2#c����_��� �C�c(\BCCFG !�[~���p!Ekem`eo���o �o�o�o�o�o�o ?*cN`��� ������;�&� _�J���n�����ˏݏ�Ȍ��ɏ*�<��� �r�]�������H�ڟ ԯ�����,��P� >�t�b�������ί�� ����:�(�J�p� ^���������ܿʿ� � �6���J�\�z� �Ϟ���ϰ������� �.�@��d�R߈�v� �ߚ߼߾������*� �N�<�r�`���� ���������$�&� 8�n�\���HϪ����� ����|�"2XF |��n���� �0fT� x�����/� ,//P/>/t/b/�/�/ �/�/�/�/��
??:? L?^?�/�?p?�?�?�? �?�? O�?$OOHO6O lOZO|O~O�O�O�O�O �O_�O2_ _B_h_V_ �_z_�_�_�_�_�_�_ �_.ooRo?jo|o�o �o�o<o�o�o�o <N`.�r�� �����&��J� 8�n�\�������ȏ�� �ڏ���4�"�D�F� X���|���hoʟܟ�� ����B�0�R�x�f� ���������ү��� ,��<�>�P���t��� ��ο�����(�� L�:�p�^ϔςϤϦ� �������ȟ*�<�Z� l�~��Ϣߐ߲����� ��� ���D�2�h�V� ��z��������
� ��.��R�@�b���v� ������������ N<r(ߊ�� ��\�8&�\Fz�$TBC�SG_GRP 2�"F� � �z 
 ?�  ���� ����5//Y/k+�~�$�d@� ��!?z	 H�BLk(z�&j$B$  C���/�(�/f�/Cz�/(=A�k(�333?&ff?7��i%A��/m?:80 k(�͎6S5f�0DHp?�=@�H0`j%K1�5j$�1D"N! �?�?�?�?;OJ�(I& �(nE�OLO^O�O�O�O��O�O_ [�H:Q	�V3.00�	�lr2d S	�*\PTTyk_*_ ��Q�I �Pt]�_ � �_�_�[~J2%�=Qo�UCFoG 'F�Y �"j�Lb�ROlwl�wo�o�j O�o�o�o�o�o =(aL^��� ������9�$� ]�H���l�����ɏ�� Ə���#��G�Y�� � d�v���2�����˟ �ܟ� �9�$�]�o� ����N�����ۯƯ� �zf6�BF�H�Z� ��~�����ؿƿ��� �2� �V�D�z�hϞ� �Ϯϰ��������
� @�.�d�R�tߚ߈߾� �����ߴ����>� `�N��r������ ����&���6�8�J� ��n������������� ��"24F|j ������� B0fT�x� ����/�,// P/>/`/�/0�/�/�/ l/�/�/???L?:? p?^?�?�?�?�?�?�? �?O O"OHOZOlO&O |O�O�O�O�O�O�O_ �O_ _2_h_V_�_z_ �_�_�_�_�_
o�_.o oRo@ovodo�o�o�o �o�o�o�o*�/B T����� ����8�J�\�� l���������ڏ��� �ʏ4�"�X�F�h��� |�����֟ğ���
� ��T�B�x�f����� ����Я�����>� ,�b�P�r�t�����6 Կ�����(��8�^� Lς�pϦϔ�������  ߾�$��H�6�X�~� �ߢ�\�n���������  ��D�2�T�z�h�� �������������
� @�.�d�R���v����� ��������*N `
�x��F�� ��$J8n ��Pb���� /"/4/F/ /j/X/z/ |/�/�/�/�/�/?�/ 0??@?f?T?�?x?�? �?�?�?�?�?�?,OO PO>OtObO�O�O�O�O �O�Ol�_._�O_ L_^_�_�_�_�_�_�_  oo$o6o�_ZoHojo lo~o�o�o�o�o�o �o2 VDfhz �������
� ,�R�@�v�d������� ��ΏЏ���<�*� `�N�����@_����ҟ |���&��6�8�J� ��n�����ȯگ������"��F�0�  l�p� p���p���$TBJOP_�GRP 2(8���  K?�p�	����*����@��@�� 0���  � � � � �p�� @l���	 ߐBL   �C�� D����<���E�A�S�<�B�$����@��?�33C�*� ��8œϞ� �2�T������;�2�t��@��?����zӌ�-�A�>�Ȇ��� �����l�>��~�a�s�;��p�A�?�ff@&?ff?�ff�ϵ�8� ��L���}�������:v,���?L~�}ѡ�DH��5�;�M�@�33`������>��|օ��8��a�`ự�	�D"�� ������`�r�|���"�9������g� v��x��נ������� ������0(V �b�����Lp�C�p�	��ſ	V3.0�	�lr2d��*�b��k�p{ �E8� EJ� �E\� En@ �E��E�� E��� E�� E��� E�h E��H E�0 E�� Eϒ�� �E�� E��x E�X F���D�  D��` E�P �E�$�0�;�G�R�^p �Ek�u�������(�� E������X 9��IR4! H%�
(z�`/r"p�v#���߱/��ESTPA�RSI d�����HR�� ABLE 1+*��J p��(�'Q �k)�'�(�(�o�w��'	�(
�(��(5p��(�(8�(K!�#RDI�/��??(?:?L?^5�4O�?�;�?�?O O2N�"S�?�� �:�O_ _)_;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo���@�O��7�i sO�O�O�OU?g?y?�?�?�8�"pbNUM [ 8������x� J K �"_CFG ,Y{s��@��IMEBF_�TT�!u��� �vV�ERI#�a�v�sR� 1-�+ 8$mp�k�� ;��o  ���,�>�P� b�t���������Ώ�� ���(�:���^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� � 2�{�V�h����������¿Կ���
��"�q_�Sq�v@�u� MI__CHAN�w �u} u�DBGLV���u�u�!x�ETHERAD ?�%���v ����x���(x�ROUT�p!WJ!*�H��?SNMASK���s>��255.��N��ߖߨ�N� OOL�OFS_DI� �BŪ�ORQCTRL .�{>Cw/&�T�J�\�n���� �����������"�4� F�X�j�z���������#PE_DETA�I����PGL_C�ONFIG 4�Yyiq��/ce�ll/$CID$/grp1��;M_q�9C�߮� ����,>P bt����� �/��:/L/^/p/ �/�/#/�/�/�/�/ ? ?�/6?H?Z?l?~?�? ?1?�?�?�?�?O O�n}�?VOhOzO�O�O �Oq���O�M��?_ _1_C_U_g_�?�_�_ �_�_�_�_t_	oo-o ?oQocouoo�o�o�o �o�o�o�o);M _q ����� ���%�7�I�[�m� ������Ǐُ��� ��!�3�E�W�i�{��� ���ß՟������ /�A�S�e�w���������ѯ����� ��User V�iew )	}}1�234567890J�\�n���������X5�	̿��0�2=� ��� �2�D�V�h�ǿٿ7�3�������� ���o�1�߾4��j� |ߎߠ߲���#���߾5Y��0�B�T�f�x��ߙ�߾6�������@��,���M�߾7�� ������������?�߾8u�:L^p������ l�Camera ;�1�0BT2BE�~��H������//�   ���f/x/�/�/�/ �/g�/�/?S/,?>? P?b?t?�?����� ?�?�?�?OO,O�/ PObOtO�?�O�O�O�O �O�O�?�7XىO>_P_ b_t_�_�_?O�_�_�_ +_oo(o:oLo^o_ �72+�_�o�o�o�o�o �_*<N�or� ����so���a �(�:�L�^�p��� �����܏� ��$� 6���7t�͏������ ��ʟܟ�� ��$�o� H�Z�l�~�����I��7 (	9�� ��$�6�H� �l�~���ۯ��ƿؿ ���ϵ�ǧ9��O� a�sυϗϩ�P����� �Ϙ��'�9�K�]�o���
	�0߼��� �������:�L�^� ߂��������� ��� ���5�G�Y�k� }���6������"��� 1CU���I+ ���������� 1C�gy�� ��h�յ;X// 1/C/U/g/�/�/�/ ��/�/�/	??-?� �![�/y?�?�?�?�? �?z/�?	OOf??OQO cOuO�O�O@?��k0O �O�O	__-_?_�?c_ u_�_�O�_�_�_�_�_ o�O��{�_Qocouo �o�o�oR_�o�o�o>o�);M_qm  i���� ����0�B�T�f�   v~���� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~��������ƿؿj�  }
`(  �p( 	 ��� B�0�f�Tϊ�xϚϜπ���������,���� ��oq߃ߕ� ����������c `�=�O�a�߅��� ������&���'�n� K�]�o����������� ����4�#5GY k�������� �1C�gy �������	/ P-/?/Q/�u/�/�/ �/�/�//(/??)? p/M?_?q?�?�?�?�/ �?�?�?6?O%O7OIO [OmO�?�O�O�O�?�O �O�O_!_3_zO�Oi_ {_�_�O�_�_�_�_�_ oR_/oAoSo�_wo�o �o�o�o�oo�o `o=Oas���o �o���8�'�9� K�]�o��������� ۏ����#�5�|�Y� k�}�ď����şן�8��B�"�@ �*��<�N��$�����+frh:\tp�gl\robot�s\lrm200�id��_mate=_��.xml
��� Ưد���� �2�D�V�F���`������� ��Ϳ߿���'�9� K�b�\ρϓϥϷ��� �������#�5�G�^� X�}ߏߡ߳������� ����1�C�Z�T�y� ������������	� �-�?�V�P�u����� ����������) ;R�Lq���� ���%7N Hm��������/!/3/E.g�Ν� $�r�<<w p� ?�E+ �/E/�/�/�/�/�/? �/?<?"?4?V?�?j? �?�?�?�?�?�?�?
O�8OF��$TPG�L_OUTPUT� 7P�P� h tE�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_��_�_oo'otEh ��=@2345678901Lo^opo�o�o �o�cF�Io�o�o�o /�o3ew���Ez}����� '���]�o������� ��O�ŏ����#�5� ͏C�k�}�������K� ]������1�C�۟ Q�y���������Y�ϯ ��	��-�?�ׯ�u� ��������Ͽg�ݿ� �)�;�M��[σϕ� �Ϲ���c�u���%� 7�I�[���iߑߣߵ� ����q����!�3�E�W���HA}c!������������@j/�.��p* ( 	  1oc�Q���u������� ��������)M; q_������ �7%GI[��?f�f &� �-�#/5//Y/k/ 9j��/�/H/�/�/�/ �/?,?�/0?b?�/N? �?�?�?�?�?>?�?O �?OLO^O8O�O�O�? |O�O�OvO __�O_ H_�O�O~_�_*_�_�_ �_�_�_ol_2oDo�_ 0ozoTofo�o�o o�o �o�o�o.@dv �o^��X��� �*���`�r���� ������ޏ<�N��&� ��2�\�6�H������ ��ڟt�Ɵ�"���F� X���@���(�z�į֯ �����j���B�T�� x���d������0��� Ϣ��>��*�tφ� 俪ϼ�VϨ��������(�:��)WGL�1.XML��o���$TPOFF_L�IM �����}�N_SV���  ����P_MON 8�S����2y��STRTCHK �9������VTCOMPAT���6��VWVAR �:��Y�� �� q�������_DEFPRO�G %��%������ISPL�AY���ޡ�INST_MSK  ��� ��INUSsER,���LCK5����QUICKMEyNY���SCREx���7�tpsc��5����ҩ��_��ST*��RA�CE_CFG U;��Y���	z��
?���HNL C2<��`� �� L^p�������
��ITEM 2�=8 �%$1�23456789y01  =<)xOai  !ow��3�z�� A//w)/��v/ ��/��/�/M/=/O/ a/{/�/�/�/U?{?�? �/�??'?9?�?]?	O /OAO�?MO�?�?�?qO �O#O�O�OYO_}O�O X_�Os_�O�_�__�_ 1_�_og_'o�_7o]o oo�_{o�_	oo�o?o �o#�oG�o�o�o Sk��;�_ q:��U��y���� ���%��I�	�m�� ?�ŏ��Ǐُ���w� !�͟��i�)����� ��+�՟�������ů A�S�e��7���[�m� ѯy����п+��O� �!υ�7ϩ�����߿ ��ϯ�����K���o� �ϓ�߷�c߉ߛ��� ��#�5�G�����}�=� O��[����߲���� 1����g�����f����S��>k��g  �k� ����
 ���������UD1:\�&��}�R_GR�P 1?� 	 @��q��m������� �  �&J5nY?�  ��� ����/�// '/]/K/�/o/�/�/�/�/�/�/	9�?%?~{�SCB 2@�� tq?�?�?�?��?�?�?�?Oq�UT�ORIAL A���LOv�V_CONFIG B�����	�O[MOUT?PUT C���@���O�O__ 1_C_U_g_y_�_�_�_ �_�_�A�O�_oo1o CoUogoyo�o�o�o�o �o�_�o	-?Q cu������o ���)�;�M�_�q� ��������ˏݏ�� �%�7�I�[�m���� ����ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������ ��'�9�K�]�o߁� �ߥ߷���������� #�5�G�Y�k�}��� ��������O�E�O'� 9�K�]�o��������� ����������#5G Yk}����� ��1CUg y������� 	/-/?/Q/c/u/�/ �/�/�/�/�/�/?/ )?;?M?_?q?�?�?�? �?�?�?�?O?%O7O IO[OmOO�O�O�O�O �O�O�O_ O3_E_W_ i_{_�_�_�_�_�_�_ �_o_/oAoSoeowo �o�o�o�o�o�o�o o+=Oas�� �������& 9�K�]�o����������ɏۏ���������0�B�,��m� �������ǟٟ��� �!�3�E�W�i���� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sτ��ϩϻ��� ������'�9�K�]� o߀ϓߥ߷������� ���#�5�G�Y�k�}� �ߡ����������� �1�C�U�g�y���� ����������	- ?Qcu����� ���);M _q������ �//%/7/I/[/m/ /��/�/�/�/�/�/ ?!?3?E?W?i?{?�;��$TX_SCR�EEN 1DD��,��}�ipnl/�0gen.htm�?�?�?�OO%O��Pa�nel setup)L}�)OjO|O�O�O�O�OXONO�O_ _1_C_U_�Oy_�O�_ �_�_�_�_�_n_�_-o ?oQocouo�o�_,o"o �o�o�o)�oM �oq�����B T��%�7�I�[��  ������Ǐُ��� t�!���E�W�i�{��������>UALRM_MSG ?�9��0 ���*�� 5�(�Y�L�}�p��������ׯʯ����ӕS�EV  ��Q�ђECFG �F�5�1  ��%@�  A�� �  Bȍ$
   ��#�5��ƿؿ��� � �2�D�V�h�v�]��GRP 2Gg�; 0�&	 �����ӐI_BBL_N�OTE Hg�T��l�"�0�!s���DEF�PROݐ%� (%�:ߖ (�a�L� ��pߩߔ��߸�������'��K���FKE�YDATA 1I<�9��p v��&�ϰ�����������,(�+��$�OI�NT  ]3�5� OOK T��{�b�NDIRECT����� CHOICE�N���F�UCHUP�����F�RE INFOOaH� l�������9 ]o ���/frh/g�ui/white�home.png�p������ } �point��*/</N/`/r///l7ook"g /�/��/�/�/�/*indirec/4?F?X?xj?|?.clos��'?�?�?�?�?O*t?ouchup$?<O�NO`OrO�O.arwrg#?�O�O�O�O_ �H#_5_G_Y_k_}_�_ _�_�_�_�_�_o�_ 1oCoUogoyo�oo�o �o�o�o�o	�o? Qcu��(�� �����;�M�_� q�������~��ӏ� ��	��-�4�Q�c�u� ������:�ϟ��� �)���;�_�q����� ����H�ݯ���%� 7�Ư[�m�������� D�ǿ����!�3�E� Կi�{ύϟϱ���R� ������/�A���S� w߉ߛ߭߿���`��� ��+�=�O���s�� ������\����� '�9�K�]��������з�����v���>����# 5WiC,U� M������ <N5rY��� ���/�&//J/ 1/n/�/g/�/�/�/�/ ���/?"?4?F?X?g� |?�?�?�?�?�?�?w? OO0OBOTOfO�?�O �O�O�O�O�OsO__ ,_>_P_b_t__�_�_ �_�_�_�_�_o(o:o Lo^opo�_�o�o�o�o �o�o �o$6HZ l~����� �� �2�D�V�h�z� �����ԏ���
� ��.�@�R�d�v���� ����П������/ <�N�`�r��������� ̯ޯ���&���J� \�n�������3�ȿڿ ����"ϱ�F�X�j� |ώϠϲ�A������� ��0߿�T�f�xߊ� �߮�=��������� ,�>���b�t���� ��K�������(�:� ��^�p����������� Y��� $6H�� l~����U��� 2DV-��X�-�������}���,�/
/�/.//R/d/ K/�/o/�/�/�/�/�/ ??�/<?#?`?r?Y? �?}?�?�?�?�?�?O �?8OJO)�nO�O�O�O �O�O��O�O_"_4_ F_X_�O|_�_�_�_�_ �_e_�_oo0oBoTo �_xo�o�o�o�o�o�o so,>Pb�o ������o� �(�:�L�^�p���� ����ʏ܏�}��$� 6�H�Z�l��������� Ɵ؟����� �2�D� V�h�z�	�����¯ԯ ������.�@�R�d� v���_O����п��� ��*�<�N�`�rτ� ��%Ϻ��������� ��8�J�\�n߀ߒ�!� �����������"�� F�X�j�|���/��� ����������B�T� f�x�������=����� ��,��Pbt ���9��� (:�^p�� ��G�� //$/ 6/�Z/l/~/�/�/�/��/���+�������/?=�/7?I?#6,5Oz?-O�? �?�?�?�?�?�?O.O ORO9OvO�OoO�O�O �O�O�O_�O*__N_ `_G_�_k_�_�_���_ �_oo&o8oG/\ono �o�o�o�o�oWo�o�o "4F�oj|� ���S���� 0�B�T��x������� ��ҏa�����,�>� P�ߏt���������Ο ��o���(�:�L�^� ퟂ�������ʯܯk�  ��$�6�H�Z�l��� ������ƿؿ�y��  �2�D�V�h����Ϟ� �����������_�.� @�R�d�v�}Ϛ߬߾� ��������*�<�N� `�r��������� �����&�8�J�\�n� ����!����������� ��4FXj|� ����� �BTfx��+ ����//�>/ P/b/t/�/�/�/9/�/ �/�/??(?�/L?^? p?�?�?�?5?�?�?�?� OO$O6O�8K}�����aO@sO�M]O�O�O�F,�_ �O�__�O2_D_+_h_ O_�_�_�_�_�_�_�_ �_oo@oRo9ovo]o �o�o�o�o�o�o�o *	�N`r��� �?�����&�8� �\�n���������E� ڏ����"�4�ÏX� j�|�������ğS�� ����0�B�џf�x� ��������O����� �,�>�P�߯t����� ����ο]����(� :�L�ۿpςϔϦϸ� ����k� ��$�6�H� Z���~ߐߢߴ����� g���� �2�D�V�h� ?������������ 
��.�@�R�d�v�� �������������� *<N`r�� �����&8 J\n���� ����"/4/F/X/ j/|/�//�/�/�/�/ �/?�/0?B?T?f?x? �??�?�?�?�?�?O O�?>OPObOtO�O�O 'O�O�O�O�O__�O :_L_^_p_�_�_�_}���[�}�����_�_�]�_o)of,Zo~oeo�o �o�o�o�o�o�o2 VhO�s�� ���
��.�@�'� d�K�����yﾏЏ� ���'_<�N�`�r� ������7�̟ޟ�� �&���J�\�n����� ��3�ȯگ����"� 4�ïX�j�|������� A�ֿ�����0Ͽ� T�f�xϊϜϮ���O� ������,�>���b� t߆ߘߪ߼�K����� ��(�:�L���p�� ������Y��� �� $�6�H���l�~����� ���������� 2 DV]�z���� ��u
.@R d������� q//*/</N/`/r/ /�/�/�/�/�/�// ?&?8?J?\?n?�/�? �?�?�?�?�?�?�?"O 4OFOXOjO|OO�O�O �O�O�O�O�O_0_B_ T_f_x_�__�_�_�_ �_�_o�_,o>oPobo to�oo�o�o�o�o�oh��{������ASe}=��sv,���}� ���$��H�/�l� ~�e�����Ə؏���� � �2��V�=�z�a� ������ԟ����
��� .�@�R�d�v����o�� ��Я�������<� N�`�r�����%���̿ ޿��ϣ�8�J�\� nπϒϤ�3������� ���"߱�F�X�j�|� �ߠ�/���������� �0��T�f�x��� ��=���������,� ��P�b�t��������� K�����(:�� ^p����G� � $6H�l ~������� / /2/D/V/�z/�/ �/�/�/�/c/�/
?? .?@?R?�/v?�?�?�? �?�?�?q?OO*O<O NO`O�?�O�O�O�O�O �OmO__&_8_J_\_ n_�O�_�_�_�_�_�_ {_o"o4oFoXojo�_ �o�o�o�o�o�o�o�o 0BTfx� �������,�@>�P�b�t���]����]������ÏՍ����	��, ��:��^�E�����{� ����ܟ�՟���6� H�/�l�S�������Ư ���ѯ� ��D�+� h�z�Y����¿Կ� ����.�@�R�d�v� ��ϬϾ�������� ��*�<�N�`�r߄�� �ߺ���������� 8�J�\�n���!�� �����������4�F� X�j�|�����/����� ������BTf x��+���� ,�Pbt� ��9���// (/�L/^/p/�/�/�/ �/���/�/ ??$?6? =/Z?l?~?�?�?�?�? U?�?�?O O2ODO�? hOzO�O�O�O�OQO�O �O
__._@_R_�Ov_ �_�_�_�_�___�_o o*o<oNo�_ro�o�o �o�o�o�omo& 8J\�o���� ��i��"�4�F� X�j��������ď֏ �w���0�B�T�f� ����������ҟ����� ���� ���!�3�E��g�y�S�,e���]�ί�� ���(��L�^�E� ��i�������ܿÿ � ���6��Z�A�~ϐ� wϴϛ������/� � 2�D�V�h�w��ߞ߰� �������߇��.�@� R�d�v������� ������*�<�N�`� r�������������� ��&8J\n� ������ �4FXj|� �����/�0/ B/T/f/x/�/�/+/�/ �/�/�/??�/>?P? b?t?�?�?'?�?�?�? �?OO(O��LO^OpO �O�O�O�?�O�O�O _ _$_6_�OZ_l_~_�_ �_�_C_�_�_�_o o 2o�_Vohozo�o�o�o �oQo�o�o
.@ �odv����M ����*�<�N�� r���������̏[��� ��&�8�J�ُn��� ������ȟڟi���� "�4�F�X��|����� ��į֯e�����0��B�T�f��$UI_�INUSER  �������  g��k�_MENHIS�T 1J���  (���?@(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1���+�=�Oπ�)��631�IE,2Pϣϵ����y*d�v�edit��?PROG,1��"�H4�F���'��v�2�����ߩ߻����� m��962��'�9�`K�]������36� �������p���
�� .�@�R�d����������������{�۱{� *<N`ru�� �����& 8J\n��� �����"/4/F/ X/j/|//�/�/�/�/ �/�/�/�/0?B?T?f? x?�??�?�?�?�?�? O��>OPObOtO�O �O�?�O�O�O�O__ �O:_L_^_p_�_�_�_ 5_�_�_�_ oo$o�_ HoZolo~o�o�o1o�o �o�o�o 2�oV hz���?�� �
��.�O+Od�v� ������������ �*�<�ˏ`�r����� ����̟[����&� 8�J�ٟn��������� ȯW�����"�4�F� X��|�������Ŀֿ e�����0�B�T�?� Q��ϜϮ�������� ��,�>�P�b���� �ߪ߼������߁�� (�:�L�^�p��ߔ�� ��������}��$�6� H�Z�l�~�������� �������� 2DV�hze���$UI�_PANEDAT�A 1L�����  	��}/frh�/gui�dev�0.stm M?�connid=0� height=�100&_� ic�e=TP&_li�nes=15&_�columns=�4� font=2�4&_page=whole� �h�?)prim/X  }[����� )���#/ 
/G/Y/@/}/d/�/�/ �/�/�/�/?�/1?h����  �   +���i�cgtp/f�lex� �?_width=� �� �2�3� 1d�oub� 2;?8ual�?�?kO.O@O ROdOvO?�O�O�O�O �O�O�O_*__N_5_�r_Y_�_�_�_�_?=  � �U�Oo$o6oHo Zolo�_�oO�o�o�o �o�ouo2D+h O������� 
���@�'�d�v��_ �_����Џ���Y� *��oN�`�r������� ��!�ޟş��&�8� �\�C�����y����� گ�ӯ�����F�X� j�|������ĿֿI� ����0�B�Tϻ�x� _ϜϮϕ��Ϲ���� ��,��P�b�I߆�m� ���/������(� :�L��p�㿔��� ������U��$��H� /�l�~�e��������� ������ DV�� �ߌ�����9 
}�.@Rdv� �����// �</#/`/r/Y/�/}/ �/�/�/�/cu&?8? J?\?n?�?�/�?�?) �?�?�?O"O4O�?XO ?O|O�OuO�O�O�O�O �O_�O0_B_)_f_M_�_�/?}��_�_�_�_
oo.o)�_So�5 Boo�o�o�o�o�o@o �o�o!W>{ b���������/��83;�$U�I_POSTYP�E  5?� 	 ;����a�QUICKME/N  p�����c�RESTORE� 1M5�  �*default�;�SINGLE~ԍPRIMԏ�mwintpe�,1,PROG,1<�p�������I��� П�������<�N� `�r����"������ ϯ��
��.�@��d� v�������O�п��� ��ï%�7�Iϻ��� �ϨϺ���o����� &�8�J���n߀ߒߤ� ��a�������Y�"�4� F�X�j������� ��y�����0�B��� ��a�s���������� ����,>Pbt��������S�CRE��?���u1sc��u2!3!4!5*!6!7!8!�wTATl�� ă<5Y�USER�ks#�3�4��5�6�7�8��a�NDO_CFG Np��P�Qa��OP_CRM5 c �U&a�PDd���No�ne���_INF�O 1O5f 0%��/�8o/�/ �/�/�/�/
??�/@? #?d?v?Y?�?�?�?�?���S!OFFSET' Rp�j!�?� ���!O3OEOWO�O{O �O�O�O�OO�O__ _J_A_S_�_w_�_�_ �Kŏ�]�_
o
�_/o>�8UFRAM%�/�P!RTOL_AB�RTSoN#kbENB�toehGRP 1S�����Cz  A��c�a��o�o�o�o�"v,>cj��U��h#!�kMSK  ��ef!�kNPa%�^)�%�_��e_EVNs`�t&�v��2T�;
 h#!�UEVs`!t�d:\event?_user\�7�#C7<�o� Fq�/��SP5�:�spo�tweldl�!�C6��r���#�t! �K�	�>��q��-� �q���Q�c�ܟ�� � ����ϟH��l��)� _�����د����˯ � �D���z�%����� [�m�濑�
ϵ�Ǻ�?WRK 2U�a#8�nπ� \ϥ� �ϒ��������#��� G�Y�4�}ߏ�j߳��� ���������1��B��g�y��$VARS�_CONFI�Vn�; FP����CMR�b2\�;xy� 	$ ��0�1: SC13?0EF2 *�	�J���X�ȸp� [ #!?�p@pup"p�z� o]�g����������h����`�uA�����,� B���G�K��l ���_����� ��2�hSe��Q����IA_�WOF�]^-˶,�		�Q;%/+'G��P �> ���R�TWINURL k?��������/�/�/�/�/�/�SIONTMOU�� ��%�^S۳�S۵@�a FR:\�#�\DATA؏  ��� UD1�66LOGC?  �\9EXh?'q' B@ ���2�{1U��?{1�?�?θ �� n6  �������2zt��`F��  =����BA��?@|=TR�AIN�?AQB�d�CpBEFF/B�0�(:��_� (��I �M��O�O�O__P_ >_t_b_|_�_�_�_�_\�_�(_GE3`�/C�
�`'p4b
g�0�RE!0a�i���L�EXdb����1-�e�/VMPHASOE  ���C ���RTD_FIL�TER 2c� �&��T��o +=Oas���� �o������1��C�U�g��)SHIF�TMENU 1d^�K
 <�<%�?ŏ2����ɏ�ُ �8��!�n�E�W�}� �������ß՟"����	LIVE/S�NA��%vsf�liv�n4��>�# SETU��W�menum�r��ѯ��"��3e`+|�M�O3ftn�z��Z�D�gQm˳<�A��P�$WAITDINEND8L!�>k�OK  �醼� :��S����TIM.5���Gr�� ��%˴��ӿ�򿆸RELE�a5��k�x�/6m�_ACTJ��4� !��_?1 h���%�5߅���R�DIS����$�XVRnaitn��$ZABC��1jNQk ,�@�2=�n�-ZIP2kQo����)���MPCF_G 1l���l!0L"��q�7�MP�m����P����؋��`�*�  ���f<�(G��3ޙ��?��6�� 168Ÿ6�ff�H�C	����	(>B���h��0�Q�����?���0B���r;T�ǯo@�S&������
�?�.�@�?m�p9��������C��@��D"(>�N���a�3�]��2��@l�PJ\r��D�)�O�4%:�\�[�(`68<�6W+�l���?��������0G��g8���a��'���J�p`n��_C_YLIND�aoR�� �p6 ,(  *o�w3l���� ��// '.iJ/�n/U/g/�/ ��/�/�///?�/�/ F?-?j?Q?�/�?�?r�Cp*� �g� �?L^���6O!OZO?Ih�?�O?G��AA�=�SPHERE 2qO�?�OT?�O_ �O:_�?�Op_�_�/�_ E_+_�_�_ o�_Y_6o Ho�_�_~o�_�o�o�o��oo�o ��ZZ�� ��