��   ��A��*SYST�EM*��V9.1�035 7/1�9/2017 �A   ����BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG����DHCP_CTR�L.  0 �7 ABLE? $�IPUS�RET�RAT�$SE�THOST��N�SS* 8�D��FACE_NU�M? $DBG_�LEVEL�OMo_NAM� !� {FT� @� �LOG_8	,CM�O>$DNLD_FILTER��SUBDIRCA�PC��8 . �4� H{ADD�RTYP�H N�GTH�����z +LSq D� $ROBOTyIG �PEER�ބ MASK�MR�U~OMGDEV|��PINFO��  $$�$TI ���RCM+8� ?$( /�QS�IZ�!S� TA�TUS_%$MA�ILSERV �$PLAN� <�$LIN<$C�LU��<$TOޥP$CC�&FR\�&YJEC|!Z%�ENB � ALkAR:!B�TP,��#,V8 S��$�VAR�)M�ONx�&���&APPL�&�PA� �%��'PO�R�Y#_�!�"AL�ERT�&i2URL� }Z3ATT�AC��0ERR_oTHROU3US�9H!�8� CH- c%�4wMAX?WS_|1w��1MOD���1I�  �1o (��1PWD  � L�A��0�ND�1T{RYFDELA-Cx�0G'AERSI���1Q'ROBICLK�_HM 0Q'� XML|+ 3SGFRMU3�T� !OUU3 G_�-COP1�F33ĿAQ'C[2�%�B_A�U�� 9 R�!U{PDb&PCOU{!��CFO 2 �
$V*W�@c%D_UMMY1TW2?��RDM* �$DIS��SN,#	3 �	o!�"�%"_WI�CTZ�_INDE�3�PO�FF� ~UR�YD���S�  
 �t Z!RT�0N�cD�bHOUU#E%Af:a"f:a1f�LOCA� #$�NS0H_HE����@I�/ 3 �$ARPH&�_IPF�W_* O�F�PQFAsD90��VHO_� 5R{bEL� P����90WORA�$ACCE� LV�O#�FS1�IC�E�3p� �$�c ? ���Rq��%
��
Gp�PS�APwo# ��cqIz0ALOaq'0 Vpx
���F�����{p�r�u�$� 2�{��]r�} �p�� �}��!YqA�����$� _FLT�R  oy�p *��������U��$�}2U��bSHA�R� 1�y P=���t���C� �g�*���N���r��� 埨�	�̟-��Q�� u�8�J���n�ϯ��� ���گ�M��q�4� ��X���|����޿� ֿ7���[��g�Bϐ� ��x��Ϝ�����!��� E���{�>ߟ�b��� ���ߪ߼����A�� e�(��L�����ﰦ��Y�z _LUA1}n�x!1.B�0���A�1R����255.��I���	��u@�2G�Y���m��������3��Y�6  ����	��47Y�@� ]o����5��Y�&�����6 'Y��M_q�����7!"��������܀ �� Q�	 ���<9/n/�/S/��/�/�/�/�/�/��P �/.?@?R??v?�?�?@�?k?�?�?�?��?����u>O)L
ZD�T Status��?MO�O�O�O��}�iRConnec�t: irc�D/?/alertkN�O _"_4_�G}Ob_t_�_P�_�_�_���sP�"��d���_�_	oo -o?oQocouo�o�o�o��o�o�s$$c96�2b37a-1a�c0-eb2a-�f1c7-8c6�eb56b02a8  (Q_"uOF�Xj|�����((�0"�r2J�u �v3C5 �,$=��� 3��%��I�0�V�� f�����Ǐُ����� !���W�>�{�b���q0!/� DM_!�/��SNTP��	��%u�����}��������#ϓUSTOM �
�����/  ���$TCPIP�����0H'%!�TKEL'�/�,!���H!T�R�����rj3_tpd�)O 4��!K�CLƯ˫���v!CRT%��l�'"���!CONS�m�̪ڡib_s'monu�i�