��  	NK�A��*SYST�EM*��V9.1�035 7/1�9/2017 �A  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ����AIO_CN�V� l� RA�C�LO�MOD�_TYP@FIR��HAL�>#INw_OU�FAC� �gINTERCEmPfBI�IZ@�!LRM_REC�O"  � AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� ."��!_�IF� P �$ENABL@�C#� P dC#U5K��!MA�B �"�
f� OG�f d �PPINFOEQ�/ �L A q?1R5/ H0�f69EQUIP� 20NAM�� ��2_OVR��$VERSI�� �!PCOUP�LE,   $�!PP_D0CES�0�!�81�!"PC�> [1	 � �$SOFT�T_�ID�2TOTAL7_EQ� $@%@�NO(BU SPI_OINDE]=EX�2SCREEN_�4��2SIG�0��?�;@PK_FI�0	$THK�Y�GPANE0D �� DUMMY1"d�D�!�E4�A!�RG1R�
 � _$TIT1d  ��� �Dd�D� �D�@��D5�F6�F7�F8
�F9�G0�GW�A�EW�A�E.W18W �F�LW1VW2aR!SB�N_CF�! 	8� !J� ; 
2f1�_CMNT�$�FLAGS]�C�HE"� � ELL�SETUP �� $HO�0 P�R<0%3cMAC{RO?bREPRHhD0D+<@�bb{jd^ UTOB U��0 9DoEVIC�CTI�0��� @13��`B�ce#VAL�#IS�P_UNI��`_�DO�f7�iFR_FZ@K%D13�A�c�C_WA�d�a+z�OFF_�0N�DELXxLF0�a�Acq��b?�adp�C?�1`yA�E�C#�s�A�TBXt���MO<� XsE � [�MXs���qREV��BIL�w19��AXI� �rR 7 � OD5`��$NO�PM@��p�
� �/�"`�� +�V�  ��X@D�T p �E RD_E
��q�$FSSB�&$CHKBD_SE�e�AG� Gj2 "_��TB��� Vxt:5p}�C �a_EDu >� � C2�eA`S8p�4%$l �tt$OP\@B�bq!�_OK��US�1P_C� !��d��U S`LACI�!�Rae���� �aCOM9M� �0$Da�w��H@dp ��O�B�IG�ALLOW� �(KD2�2e@VA�Rݕd!PAB =m��BL#@S � ,�K�a��`S+p"@M�_O]"���C�CGXpN�!o $��_ID�L�`��$�� B��)AS� c�CCBD	D�!{�I����LPz�|84_ CCSCH�1�` OOL��`�M�M��S�C�s$MEA�P\t�`Tg`�!���TRQ�a�CN����FS3k��!/0_F��( )��p���U� �!B �CFn�T X0GR�0���M�qNFLIx�u�@UIRE�x���!� SWIT=$�(�N'`S�"CF_��G� �A0WOARNM pP���r�PLX��NST� �COR-���`FL{TRܵTRAT �TR�� $ACC�a�� �r$OcRI�.&��RTj`�_SFg CHG*x@I��Tp�A
�IF�T�!���>� � �#a����HDh�Rq��2B�BJ; �C����3��U4��5��6��7��e8��9�!h�CO�S <� i�{���x3�2-�LLEC��}�rMULTIr�
2ʓyA
2FS��I�LD	�
1v�B@T_��R  4� S�TY2pbܖ=�)�2ܐ��`��0� |A06$��`@�ޔa`�* ��TOx�:�E,�EXTB�e�p?��Be�f22n0,����0��R�.'�������� �"�/%9a9�����cg����� ���A�C�?�ME� �� q�Ջ��! L0���� ��cpA��$JOB�Ȱ�l�K�;IG��" d{�^� p�����-'��8�嗷��ACO_M��b#� t{�F� �CNG�AiBA� w�DɁ M
/1Bk�j0W�F@�yP�`zm÷$ϰ$��t�a�"��
2J"�_R�a"C��J%���J�D/5CԽ��Fn@b �W�P�O�л!% \0RO�6i(��S��O_NOM_ �`n#�jc�Aᦰ������ T0�&"�@<�U��Pk��e�RA@@n �3"��?�
$TF�<�D%3S�TP�pU�1���%�%�H�b�T1Y*E������#��p�%���A�YNT�"�TDBGDE�!'���PU�@��=�82C�AX�㟲[uwTAI�cBUF��8+ѳ!\1( ����&��PIӄ'�P�D7MC8MP9� S6F>D7SIMQS�@�wKEE�3PAT ���"�"#�"m�A�Cb%)���pw`JB��U�vaDEC�:[�58*�A�$* �����v�MP��$G- �G��_e jc��1_�FP�e TCJFS W�MEb��_D?#� J��V��V��Q��FJR�F�V�SEGFRA�6�O����@T_LsIN���CPVF�q;��`t �$+G�l��B�����B"r�2�,` +,��ܵQ�� F�P�0'`�bRTm�aY�1SIZ��r�}T\V�TgS- �Z�YQRSINF� ІC�@�@�I�\�@�Xk@�@Le�8d )@fCRC��?sCC�e�@6hJA�� JBۢqdeJA�Hh�Q"eD����|iC�kcp���~D�`���f< �hE�V�f�F�a_}EFo@Nv�@�1ܶ�h+�,݀�C%�+d!V'SCA��e Ajv��Rɰ1�C�-��	��MARGh�C&�F�@6�_AD�Q��_@LI����kb`���8J|��#`r�.� <�Nߌ�S�t5��� �HANCq�$LG��O���{�4 ��B(�A�< ��0R�rrC~�ME�1���)0fy�RA��~�AZ��ň�`@%Oa�FCT h��p)���eb_@�0� ADI�O���A ��<X������L�S���B�BMP��D�PY�7A4�AE�S�P�cB H�U�0M�MENU�/��T#IT�q���%��AH�!)1��L�Ѐ�0d,�Q��OR	R$����	P  ��Ou���O��4%�������E�V/#(У DBPX�WO�P��1)�$CSK�2���T9�wTRL�2 �� �AC�@A�&�IND&� DJ8��_kp1���;���PL	Q��2WA��ΠE(�D��!ۧ�!�R���UOMMY9"��1�Л �DBρ�3�c�)1PR�Q 
p�������4 �ж'$��$�Q �L<�5I�[�c���6o����PCr�7����ENE���q8����R�ECOR��9H�&�C#� 4$L��5$<�2���0�@���A�_DJ�?0ROS� 2��{�m�`�Iñ�;�a�PA/�|��BETURN_gcMR��U� ��C]R.�EWM�B�0�GNAL� 2$L�A]�Ş6$P���7$P���8���!M`C�Đ��DO�@��)��Kb/ƟGO_AW��@�M�Oޑ:���u�CS�S_CN��Y��:`Y��T@��Z�ID'���2]�2k�N�Oд�D��`I:� �; P $��R�BoR�PIk�PO��I_BY!�����yT�RD�HNDG��< <�A��c@<�SO DSBL��S��6�l���F�LS�q=� H��060k�TO3FBm�$FE9��砒�l�Dө�q>b�D1O7A,S`�MC@��[��4��⚒H�W�( �MY7��SLkAV�r?�BIN� ���63�֭�_�@P!P�`@���А�� А�u��!��Z�?�BY�I$����W��΀�NTV3[�VE4�SKI��A�$�3��2�B7AJv7A��~DSAF�ZE�_SV.�EXCL�U�� �rONLD��>Y��]��EA��HI_VI���PP+LYӠR�sH\0Q��l_M$"��VR�FY_��jM�s�$IO�0��#`1��B���O��oLS(p����4�!�l�)�@�PK�$J��?AUTOCN� ���4l���[WCHD�\�5�_����AF&9�CP��TT�!�8=�6�j� AӰf�r\!_@w  s����SGp B �* CUR����1 � �� �@��F��F�>�ANNUN��= #l�������d��1).!#`6*R&�EF��I��C @�F"Ŕ`OT�����@����n M��NIC�DT��",W� �AU��$DAY�L�OAD����"�5��#EFF_AXIJ\�EӰ�Q��O0|����_RTRQ�q�F DWq�H0�R�T3@\45 2Ep�@�wC1�� �A�p�81�qG 0K!�1A0�T�2�/�DU��/�]�|�CAB�qH|"��p@�0P@ID�@P�W�s�5@Q_@V��V�_�0z0Ҁ�DIA�G��qI� /$V��YUT�GHA�Q��NJ��RRʲ�!�T�VE� SW��A���P�0�BC5z0F��PC1OHY5�1PPL�@ cIR���RB�P��2�3�q�� aL �BBAS;�G��Ҁ�E�ք�5z0H�H0J��UR7QDW�EMS�@HU�AKp�EsB�TLIFAEkpT#rP�~RN�Q b�U.!�SbZq��."�C��3�N��Y��p��FLAh�/ O�VJ��VHE��BSOUPPO����~Rb��_�T��Q_Xw�(d.�)gZ&jW&j��`)g�.!'�.�XZ���3��QY2�hC �TF�G�MEN�pKD8�@��?�J `��CA�CHE%w�bSIZдV�PH��N��UFFI%`Z�kt��2�6"�8�MSW�eK 8�KEYoIMAG��TM!�@��Kq��Fv��t��OCVIE�@�L � �L���w�?� 	�6��M�P0��ST��! �r堻t�t0�t0>�pEMAILp�\�x�!��qFAUL�"qN�rZÖ�COU��䃐�T�2AO<' $&���S�0�0;IT��BUF�gw�P�g��Ӑɐ�PBR����Cv�A�'���4�SAV��_�d@�bw�F���'�2&P�����D�5�_R���� ��OTN�V�3P� ����( �n�h�F� XR�C�у_G�S
u�YN)_�A5pP�2D�ճ�����BM�2�PTz�F���E��H(���4qQ�` Gs��!&�+���s�����4qR������C_E���KU���� ��RCq����D�SP[v�PCF�I�M��=�c�x�<@U`��PTř �pIP��d��ADߐ=�TH�ȋ�0�#0TH�=�HS{DI:�ABSC���`ɰVM����#�,�34NV*G��H�`:�R�F�Aj�d���G���SC.B�����MERe�FBC�MPe�ET� �S9rFU`DU`F�p��vb0CD3�ؽ�����o�NO44qTP0��޲�%�ܴ�%PS۵Cߐ�C7!�1ٳ'��5pUH *�L R����&�h�P W�� ^Ė\Ʈ!\�1\�1�\�#q\�7Y�8Y�9PYʅP[�e�1r�1�U1��1��1��1��U1��1��2��2e˪r�2�2��2��2���2��2��2��3J��3e�3r��3��U3��3��3��3��e3��4��XT?A4qV <�������V���VŌ��� �����FDR.DWT2�V�~R���.~RREMg@Fq��B�OVM��A�T7ROV�DT��4�MXC�IN��P3�N+AINDR��R
~�<ޠj�$DGR��C�=�p�UtADX6=�R�IV��R�BGEA-R�IOkEK�TN����1iXa gp`>�SZ_MCMy`~Q� �F�PUR��X� ,�u�? ��Pz?P �A?PE� X�q��t�R��Y� 3PP:�;@�RIµ�_�ETUP2_ Z 0^�TD�����hp��l�_�BACv�G[ T�p_�ɔ)Ú�%�#!à��IFI��A��t�E��@PT��BߑFLUI�d�\ � ��w(�UR  Q���R����U�CC�h0I��$�S@k?x�JƐCO���VRT��� x$�SHOg1= �AS�SΠ��U����BG_�����������¬�JDATAZ2A]�FU;1���5$2ەJ�`2A^ �|��NAV*�)���� �S�r�S?$VISI��SC*�SEv ��5UV� O�1/1B'xe=@�&$PO� �I�A�FMR}2��_ �� Ͱ�2��א�&�����+���U�_����h@IT_:��f@�M������DGCL�F�EDGDY�8L	Dh��5�V���Tְ�� �e`+�O9 �T�FS���ta �P��+Bדj�$E#X_+ABH+A1F�9���R,@3dK5dF�G���%b �` ��S�W��O9VDEBU1G��A	�GR� ��U[�BKUf�O1n.� �0PO30��I�@���E�@M�L�OO:�QSM_0E⬂��p�P_E �c x@!rpT�ERM4Ud=U�AO�RI��9Pe=U���SM_Đ�9P�f=U��* |Xg=U���?�UP}rhg� -o�2c��KS�Pd� G�Z�0E�LTO�q$US=Es�NFIG�b�Q�; �A��bT�Te$U;FRʒ$߰�Q�&`��j0OT3g"�TqA͠��EcNST���PAT¡�`[bPTHJ��E�pԂ���RARTŀ�U�Ł��r�QREL�ja�S�HFT���Qaa�h_��R����zV �P$�W�`g�1��x�a��SHI�`�4U� ��AYLO��Z�p��My �aaV!󵿠ERVd�,q��h��Ag����b�,�u�,RyCx�ASYM�����QWJg���E ��a�y���U�t�� p��e�0{v�ePv�Ip�&�vOR��M�# �@#Q�$i1"�B	V0`` `Y���HO�D�j �Gb0� ͰO�C�Q�A!$�OP�$F�J��H ��� �R:�fa�OU�acer�R_e�Ɉ�a�e$7PWR��IM�]rR_���d� {Ptc�QCUD�m�y���k� �$Hȕ!n�AD+DR��H&QGcb���|�u�-�R�"Al H��Sa��!㴕�0��ô���SES1�#�  HS���#m $� ��_D���@�^��PRM_f"F_HTTP_ްHAwn (�OBJ� lu��$��LERc�/�� o � \�痡AB_�TS⃢Sm��\KRL~$�HITCOU� ����!ƀ������ƀ.ǀSS��W�J�QUERY_FL�A�Qh�W���QAp����INCPUxB�!O2���d�I�ʔ�J�ؔJ���T�IO�LN�q��k0Cޥ!$SL�"$�INPUT_)Q�$䀙�P�# �u�SLA�1 r����ѵʹ�s���r�FIO�F_AS:Bs� $LW��aN�UzP�`ae0���@��.pHY��P��)�.Q�UOPEt `�n���b�@�b�GƘ���P��䀎ǲ� Gƿ¨��� M�qRgu lJ@sTADr^�A�TI���:��30ի`PS�BU30IDW0���7�Ԁ`6Մ���2�S`vȲ"��#���N��30>���IRCA���� w � ��1�Y��EA8��џ! ��b��ׇR{`�q<9��DAY_?�:�NTVAaN�&���8e2�&�SCA>p&�#CL��?���?Ҝ �RxjߋԀb�ա�N_��C2��?��SyȲ( �����R�?��6���(! 2x� ���Rz��R��LABSa+�301��UNI4�ePI�TY��������UJ]R�%{ ���FU@�
w�g��Ds�$�J7��O�r$J�8��7d@����7�0���8����APHMI� Q����D-@�J7J8� L_�KE\�  ��KK�LM�� | <ʰXR�?��?WATCH_� Fs\��ELD	yGL3E} f0IaVRp�֓CTR�c���BGLGO~�[ !��LG�Zw��@�@���FD�I��Q��6P �� ���@�� ��6P��p�E�P�!_CM7c�T@��A1F�q��� �(��b��@ ���'I�(`P�6P�� RSV �p`  (�@LN���"z����@TAҲ" t!��U��!m��L�#�"DAU�%E�A �4 ���"� GH������BOO����� C/�4�IaT��$�0+�RE���8SCR���0�D�I*�S `�0RGI )R�0=;��#ï�f2¤�Sc��WD4��$�#�JGM�7MNC�H��FN)�6Kn�7PRG�9UF�8�p�8FWD�8HL.ISTP�:V�8ePX�8� �8RS@IH#��; �CtC�r#�Q�x7�IU��4w7��5ȩ 8��2G�9�`PO��G#J35C��4OC�U�HRGEX�TUI�5I<����< �dQQ�3[S�0\��`?���	[�%5�`$1NO�TVANA��R=�A�I1�|�l�uDCS�༓�Sʓ�RO�XO"�WS��b�XS h[8IGN� ?��1�����TDEVzGLLB�q� c L����� m�T�$�d�:�h�w�CAd��� �����E�'���@1*�e2�e3�a�Q�P��� ����b�T��5��7�Q���@X6��;vST��R� �Y6��P^p �$ElvCl{���{vp�v��T��� L,� >���S�5�SǶ���8��EN �8�
�}2$3_ �	�i�%�X�%0� �MCu"�� ���CLDP|���UTRQLIU�p�S��Q�?�FLGgr?� �s�j�D�s���LDs�]�s�ORG0��vB���RE0����҄ʓ҄ؒ0� �� � 	\�wEN�Fs�SVe Q�, 	����,�4�RCLMCB�ҏ�T�o�4����M���� �@ $DEBUG�����T�P-�E��T�gq/�ISCv�� Yd~!qRQ, 	��DSTBO0F� ��D1	�AX�R. ��%�EXCES���l!ߒM����� ���T �ߒSCp #�*��� �_��������#�5�/�K��C \,���O0��B��LIC�tB0QU�IRE�CMO�OP����p���L�pM�� �0�<��ݣ�R��
�MND�!� �|"s"��{�D��$INAU9T51�$RSM���,`Ngro�Ca����g�PSTL�� �4��LOCvRI�>@uEX��ANGx�R����ODAQ�Ő�-��MF �B�8y�r�@�uhŜp ��SUP�uW�F�X��IGG1 � �	��soV��r�F�tb  %\s��_p ��_p�ư��C�g�᤬���`I��7� t0�MD-�K�A);��PF�Y�C�H�̳�F�DIU�F�AN�SWj1FԵa,QF�D��#)s�Ou�*�� �[ d�CU� V��Xu�����MO]1_���� ���s:Ö�&/����P��K@4#p��P��KE�B_ ��-$B����pN�D2�[G�2_T=X�tXTRA�Ss�m��<�LO� � ��b�������y�p�ҩ��r�RR2v���0 #��!A�1� d$CALII2�pG�Q��2�`�RIN���<$R���SW0`�#�m�A;BCA�D_JY���\��:�_J3N�
H�G1SP� ����PH�Bo�3n��Ѿp�����Jm����)�OvaIyMm�4�CSKP`��������J�!4�Q������_A1Z0���@EL[a���OCMP�5�PqƇ RTʑk��1�����2p1��|P�
Z�SMGZ@�2�;JG�SCLE��SPH_`4����_�����RTER|"�����INACp����^2��Y�p_N���@8=q4���5}��B�DIV5�_C�D�HE�u����`$aV�����|Q$�  �́�`�_������H �$BE�LQ ���_ACC�EL�Q�m��IORC_R�L�ŀ�NTPq<s$PS�D�Lr�N $$Y� '�!�P&>��['D�['3*"��H�_�a �� �!/��C? ��_MGoQ$DDx�! 42$FW�����%���(DE��+PPABN2'RO� EE�"�a?Q���a�����r�$OUSE_���SP���C�@�SY0�/� �qYN�A�y6���]�y1M�����R� O9LK#�4INC�����"�$	��7��
�ENCS�����"!�� INDrI*"E ��NTVE�0��+B�23_U���=CLOWLa�@��Q��5]FD�@�����p��5��C($FMOS�9`���В!t23�PE_RCH  zCO]� �G��C��`B2����f^c5i 	`��A*"UL�T����%Ep��`J[VvFTRKAqAY��S���Q*"��U�S�q���2QpMOM��	���Ȁ������#���S]#�b�D�U���"S_BCKLSH_C*"e�� �F]��3��;d�2Fj�1CLAL�`#Bő8�PpxeCHKQ�!uS�0RTY��8�D��u���_Ws�D_U	M���fC���!��cn$0LMTk�_L̀Y�dm�wE}"p{  p%u(��%Rct& XPC�A XH�p���%�eCP�z��`�'C�N_ �N`��vm�S	F��IVc2�aG�p�q*"��xCAT�nSH]� ��$�6��a�F��+!�� � PAL�d�2_P�e�S_����`�V�@��S���eJaG!�[���K@OG�w>�RTORQUU0�� �C�Y� ࢦB�Q� �_W�U�T��8���7��7�I?�IM�I�F'�*����� �VC�0�����1ೞW�ǟ���JRK�ל��떷�DB� Mt�ӷ�M��_DL�6RGRV>�7��7���H_���^ e��COSr�s r�LN ����ڕ������ �� i�Ӫ�����Z���F�MY���~�@ᆫ�2�THET0fEN�K23�\����C�Ba�CB�C��AS����i������a��SB���l�GTS��$1Cr���}��<�У$DU�`?W�����1������QQ���ws�QNE��y�I����c}	M$P�A�T�}ņ�d�o�o�LP!Hr�[�5E[�Sڕ�� ����Х[�ߦ�������V��V�ȑ��V���V��V��V��V*��V�V�H��A֠�Ҷ�;�����H��H���H��H�H�OJ��O��OJ��O��UO��O��O��O��O�O��F[���������SPBAL�ANCE��qLE6ɰH_T�SP���5���5�ЦPFUL�C9�`�H�`�Х"1=�mUTO_�`ȅ�T1T2���2N �a�-@����Qb�@�(1"��QTLPOV �>(�INSEG�A�REV��@ADI�FuUG1�,s1�*@OB"haA��W�2�-@�a �LCHgWAR2�AB��~�U$MECH���!��1��fAX�QP�Ft�vǂ�� 
p���EROB�@�CR$R��r���DO_DAT�?� < �0��O1�by1s�BE'$ON!CD_d@y0���0`u` �� %�0T@A�a�T#x2L�@�`CK�x2� CT1  %�`�N�@��8�@R3`y1������ MP�3E5 $IR���1�`8�/PN2MAI��14�2%_]#/ t!�0R,�COD7{FU�0FLAGx2ID_O`V% ��G_SUFFi� C�0�1 �1��DO� �O�(GR]��$��$��%���%��$  2u�&HV _FI-�9
3ORDA � �MMY3�6Jr2q!�$Z;DT]%�  cߟ4 *.L_�NAM�d2�DEF_It8d2��4�ST��P��0�3��5�ISD��` 0S���3�~4�E)34�q]r�2D��(b)D7D��O�/LOCKEn��#�`���1�"� UM�% d2�$�3�$�5�$B�" �C�%�3�$�4�"Q��5 �D�1�#� ���%d2�%@�3�#�G:U�(gPT  �4w�1Y��WuHtU6C	P0TE_Q�� �ZRULOM�B_�R�W0�BVI]S��ITY�BA��9O�QFRI���SFU SI�1�QE�R���W��W3�Bn�$�W�XW�[(��V��_�Ei�!EAS._cS�Á�A �GT7� 7h �TEW F�7ZuCOEFF_AO���d�\ GF�hcSU ���b�.x�$�`��C�- �cGRD� � �� $@��9XvTM^GtkE�sC,,|BER  TTDS4n0�  ��LL�$̮��ASV.D~x$ėV0��}d0� =rSETU�2c|2 � � �p6� "@ID�r��qCA�vi2�CA_A	@D�b'a�"���<@
A;@"�2�W �. R�0�qP1S�K_��c� P�&T1_USER���Yt�o �t���VEL�t�o ������I=0���MTgC|��k��  ��4 O�NORES�Jۂ�p ʂ� �4"��r�R"�XY�Z�#����DEBUz����_ERRC� ,�PpeF �c�7�Q`����`BUFINDX��P��wMOR�d� H&CU7�L���'!<1x�� 1$� r���1���2��3�G�b� � ?$SIMUL+`F �	x�VO�H�O�BJES��ADJ1U�b���AY�0��D%�OU0���\r!2=��T��pT���S�DIRX��`�/ =��`DYNH7b��T�y�R�Q�wAw��OPWO}R^� �,�`�SYSBUm��SCOPޡZ��q�U�b/ P@���PAw���q���OP� U�w�T+!A@�IMAGJ�&C��23IM��f�INE`7�~e�RGOVRD�� �x�B�PD�d��`S�P*P/C���Li@B4�|��qPMC_EE0Z�ANm�M�!A*2c19 A�P��SLS��k�� �� OVSuLSiRDEXAD�0&�2���a_�� >�� ��>�� H�]�X��b}�C� f0��Z�8Ĺsj�� @�����OH0RI�� ����* ������ɐP�L�  $�FREEȂEıR��1�Lj����yT� h ATUS�p$TRC_T|�i�@�BpJ�3��tCp A�E0k�� D& @�)�=Ҧ��>�1�`J���XED��u�Ҭ��wԳð��r�C�UP�@�1PX�j�=��D3�s��PG�ȅ�֠$SUB�2���A2���JMP�WAIT��M�J�L�OW
���$R�CVF"!��M�RXq�ɀ�CC��R������IGNR_P�L��DBTBh P��1�BWB ���UY��IG'����� OTNLN����R���dB�PN� �PEE�D��/�HADOWh ���E.�>�=���0SP�� � L&� �1^�
�l�UNIE�n�y���R��З�LY:0��<�ҿ�P��j��>�$��D��L��NPAR@T���*����P�k���bARS�IZG$0 3�1�O�� �ORMATT�¡��S��MEM2�(��UX͠���0�PL[ Ʉ� $�Ӂ^QSWITCH���aW�AS���ȑQaPLB AL_� �y i�OPBԱ�PC�D�qP���J3D�� T�`PDCKͰ�2��CO_J3 PH��BE��a��� ��b��˰ �� ��PAYLOYA�S_1Z2Z� J3AR��yfx�u��TIA4�u5�6�MOM @�����ŀBa��AD�����PUB��R�!%�!%���lg��` I$PI���U���_Xr*��]Zr*I
+I�+I�#�VA�& ��&������8}���"�HIG�"� b�[�6[�b��q�6�K3$8��39��b�SAMP�Њ��47�3b�'MOVU���,��1 ��@���4 ��6[�g �9u��������5RaN2�5INLR`k3H 9KDb�J_H6D_KK/GAMMESF��$GET}�f��iDC��
�aIB�b:�I'�$HI�TaALР��FE��X�P�L�PVLW�M<V3\�Y`VV�b�&��C���CHK���� ��I_j0.a���T QaE�W���&�Y�� �$� �1���I�pRCH�_D~���Ѓ�HpL�E������Uh?`���MSWFL��M.�SCR��7?��f��!�e �L$SVt�Pxpm��g�a�w{p�SAV��t�e/�NOCC��0�D�`�D S}![ᡑ)[� [z@K{� �%�xuD3� y0�B��6�7�2��8 �6�K8�w�u�s�1�0�T�L4`g�� � �SYLq#V�G��SU�����>��� *�V��SJ�V�q��`�� �Wp����A ��d�� �M̐��CL��������h1 �M M��aU"� � $5�Ѵ$W����P� T������"��) ��������A�@ųJX@X��O*WAZ���M ��� ��QOM�S]0BTfx�CONHb��h:C_s� |��� �`�H��H���`� u�`����E��L!,�J�b���z,�P��PMW�QU�0 �� 8��QCO�U�Q0QTH��H�O7��HYS/ ES�1�UEޠ�b�]O ��  { P܀��E��UNE�j�
8 �2u � Py�=�����a���ROGR)AX�I�2��O��<��ITK`�� �INFO��� {p����I�ȼaOI��� =(ԀSLEQ��۱��%۰s�j OS_E9DO�u � �����K�1��QEPN9U+�%�AUT
q(�COPY�10I� �pM�ANS�W˚VP�RUT� Z�NF:E�U�$GA������R� ~�� � � |����<�?USR_TS8���{TP��KLNA�4�CL��%�T�P$�OPTION��Gt�>��"R�R�S�h�R����LD@��� �� @|��A���z���M�ēPAS���P���PRG_�(Ҟю�6���= ��e�  2�PI���CH� ������/�!��_OV�bq/����M��P�T1T�W�STA�TU#I����AP|� ��MO_WA�D���X����S�P0��w��P�CR�C�� �aS��]�p��T�f��x������ M,��HEp"6�Ai��h!U k��� 1�� ��KTܥ� �< N�TRImE#SEݠNC�� a�j�Q�BѠ	�(N���Q�������G��LU��PRIp������WRK��o� ��SV����ܢ�&S2����E�XEC��R鰌� '�t�@1����(�:� '�T �� ƠELE��2� ��GA�DJ�� h9�X��MI=c������W�P�c`�3� �R�EXT_CYC�*�GN��$�9�,���LGO�S��NYQ_Fu 8"W�j@�V����C`aLA Kc��������@����PIF�!{�$��_!GKc���2�Mk��2��q!W`�LAST�!�qb��� ��z�ENAB*��EASIX!�r�2��P� G"��ay&z�@�@��S��!����Zc�"AIBCѤpE��"0V;!�&BASq�&�B]�qU@0�@p$�!~�'RMS_TR�#0WAH`3z�SP��4!��$ ��d��:7�	�� ECg� 3Dk62j792ۀ�pn�p2�7��MfDOU2�Cd��bPR�mў�GRID��C�B�ARS�&��Y#��OTO���һ`.���"'�!+BO��i�� ���L#0��Rp��<A�YESRV(��)ZDRFDIpT_ � t@�D�`�G� �G�Ъ�G5�I6�I7�I8>rAPE�PF��m��+�$VALU��#�ek$���Ai�A���U$q}�$C*��h|�AN�cR !��<�Q�qTOTA�#,� vRPW}I�1�TREGEN�Z�R���X8Q�t庡@V٠T1R�#"�Q_S�`�W�P�#V��b��!E #�0���r<�?�RS7V_H�0DAٓ`�P`S_Yqz��S��ARِ2� 
��IK�E��PRB0%�_@�+dhD�A�5փ 4��?�&�[�hSsLG�`�� @\�@P����݂6� Sy�1$DEqAUO�2�����`TEr�m��# !�Q���J�fQ�=C�IL_M�~p1V�"|Л�TQ٠�Ӥ��0C��m�V�{CF�}P_}p� �sM�y[V1�zV1�{2�{U2�{3�{3�{4�{4�zo�� o2o�w�s���p2IN��VIB�逳t��2��2��2���3��3��4��4�����r��Sf�����D $MC_9F��|	���x�fSM����7�+�F�3 9��5q� �KEEP_HNA�DD$�!f�� p�C��(���A%�����Oҡe���#�`�������RE|�r��!P��ÕڑߘU$�e���HPWD  �f�SB��+@COLLABt9PpgQ�	����O�r��N3{�\�$FLj0>�!$SYN�t��M;0C�b��PUP�_DLY��+�DGELA��!{�Y�p�ADRa� �QSwKIPe�� ���>�ORf�|��1Р�RRg��o�j2�� ��w������� �@��@��@��@�=9'�J2RG�-��bEX� T���ITS��;�b����a�b���RDCKQh��� ��R-1TOR��pp1R����!0< �m4RGEA�R û2FLG���W�L�m4SPCĲ�嵰�ds2TH2N0������� ���0POS11W�� lW���)r��U#J�[AT��CH�UjTns��IN����m4���TO�o2HOMQE��^��2����`�������� � ��3���#�5�G�Y�k߮}� ���4��†߲��������ߏ�5����/�A�S�e�w�S 氚�6����@����������7���)�;�M�_�q� +��8����� ���������S*��� � -0�óPJ��̡ڒEh��`0Y��lV�IOaq�	�IO P��R��WE��� � s�ӱu�EfT �n�$DSB��;"�eS��C��Q��S2;32�� ���y��5pICEU�"澠PE��i!PARsITRadQOPBR��h"FLOW�`TR`k qR��0i!CU�=Mh#UXTA+�i!�INTERFAC�l"_ DCHSq� tW� �00̪aT�$� 1`OM$j`sA/�<0I$�� �0An�� T� aCS �X��5(#[pEFA8�p^�[�RSP�Sq���Zp$U�SAw��q"	�EXF�IO��: �PY�%�&_�r9Q� �&WR,�7I
�0�(�M?FRIENDM1<�$UFRAM�d�0TOOL$6MY�H �2LENGT_H_VTE
4I�q<M3�0$SE:[9_UFINVQ@S����RG�2�0ITI�T7X|�e7�6G2�'G1A��#��2�7�`_2o�O_�jK <�=1�p'�>�Ce#ju��Cn�b2�1&FG �G&��Sq�r �j5�J�(�c��b����g$�wX  E_MY CT�#Hа�(����$e#Gn�W� �G��B�DDĠLOCK��E���a�AT0�=$?F 2�W��!���)1�(�2�+2
O[3�+3�*?Y�Q�)�]Y�QM� c� cVBp���U@�b1>ABTp����(S*� z�F�"k@2c�A�5�E��Nba3�}1`4ACdiPRϰgf}E��SS@���P��x�e"M� 0�0D�F4Pﲰ�T4P�W�Pe �0��
�eS��/� �	aR3!`r~�q$RUNN� SAX�@A0LH1���rTHIC�!�Ӡ4%�FEREN�auIF��#qaI�'gsM�`G1�h��tL �y�u��v_�JF�wPR@���RV_DATA�G� ��̐�� ���AL� u��v� ����q  2�� �S�O�	O� �$Ű��s��GROUǱ7�TO�Tt7�DSPN�J�OGLI�y0E_	P���O.q��� @z�K. _MIRj�d���0M�B��AP�A�iAE� ˀ5$t�SY�S���t�PG��B�RKB4&��AXI]  ��#�9��`A:�C���BSO�CB�� N>�DUM�MY160�$S}VU�DE_OP��SFSPD_OV)R�`�p1�Dy�|��OR��/ N% ��F�Nq��g�OVj�SF��p���BFٖ���p�3�.1�LCH��>��RECOVx�� �g�W��Mg�/�j�R�O�J�v�_pps @Y0VER�`.� OFS�0C�p3WD��+���J��"ą�d�TR��аE�_FDOĆMB_�CMǱ��BZ�BL b��Ѣa�dVBA�R�  O`���Gҧ�A�M�Š `�R�-�_�M頷P��_�T$SCA]�P�D�d��HBK$!3&y�IO��%����APPA |���������8��_�?DVC_DB�3�@4!�;����1	��R��3	�X�ATIEO����x�U�#\��CABs��"�3@�@<�i@��Qg�_�~3&SUBCPU��t�SR@	����% �S���S���~�$HW_C�S��%S�A�1�p�$UNI�T���ATT�RIӀ"�t�CYC=L�NECANµ��FLTR_2_F�It3T�%�QLPx��_p^p_SCTCF_�F_ܡ�*��FS$��CHA��!�������RS�D\� +�>s��� _T�PRO:����KEMe _G��T�Ҏ�Q ���QU�D�I� 5$RAILAiC��YBM �LO.�@3V��aJaX�SaX�VR�PR�S(A�`���Cݱ_	Q�FUsNC}�`bRING@`Q!j���RA��B d�	� r�	�gWAR�se�BL"A��:�� 5�/�6�/�D�A�
�t�:�3�LD@ l��A��q�Ja���TIRb��2��p�$h RIA�.AF��Pv��J���p\PR��p�MOI���DF_F0�!!��LM��FAY0HR�DY�$ORG��H��A!|�;MULCSEF0Ӄ���QV��J��J������FAN_ALMLV��WRN�HAR�D� $&�@@@��2���/��_&�3&A�U�R�ԸTO_SBR߲$[�/��߳��GMPINF�p$�Z��eRE�G�&NV" �#�D�A10��FL��}��$Ml�_u�R��p������t�"��� �0
1$�!�$Z�1���#��o� �؃EGR`7�l�'!ARI�]�T��2��6%`��AXE�Q�ROBN�RED�N�W�1�_�-0�S�Y	�a!��&S�'W�RIY0:&��STRPM�%���E��p$C$�a@B� ^�r�&5��>�OTOu9�pJ�ARYN�020��>��q�FI�?$LINK*$qJP1�Q_�#^�B%96^�x1XYZ��:�7�6OFFf�O2�w2k840BL���`�4;�5����3FI=Р�7�ao�d���f�_Jy��r��\3�A� 42;8^��ATB&Ay2^BCd�ԆDU|�A&]9��TUR� X��E>1UX� l�FGFL�P�m�4 �@�5�)�3�`� t� 1�J�pKs�M��T�3�Q���Rb�ǎ�ORQ 2�[���H]�K`뀚p�, SaeUӃY��zTOVE�Q'rM�Йq� �U#�U"�V� �X� �WИT�u������(q �Q���P
q�U�Q�W`$e#$e�S[�ERx�
�	��E� ����bd	Aa�p�5�-�<7{�x�{�AX;��r{� )���Q2�e]��i��i 0�j 0�j�0�j�0�jW@�j�@�j1�@�fg  �ig �ig �ig �ig  yg yg $yg 4yg xDyaqUyDEBU��$���U��{�s2CAB{�y���{SVn��� 
 ��<aH� ��T���T�1T� 1T� �1T��1T�WAT��A��pc@���R�3LAB�2qFU���GROg�4FB�W�B_;�If �$���0,��1�GU-�9�ANDP��Wd X�|5Zav� W�a�{1��l�Z�{0NT8� /���VELA��T�Ƒy�Ζ�$��AS�S  ���4��mPmP �k�sSIL ������Ie�|����AAVM� K �2 0�� 0  �5���g�s�d��� ��	����ͯmPB1������ߦ���� �(���.�c�u�}�A�sBStQ  1�� <Q� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�� ������������� "�4�F�X�j�|��������������ݐ$ g ������  d���IN����PR_E_EXEC �&T��0�A�IOgCNVEB ��Pk]@����IO�_p  1N�P $>����2��1�?������ $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Խ���LARMRECOV Z��&��LMDG ҷ� ��,�_IF ����� �ϥϷ���o��������/�, 
  /�X����~ߐߢߴ����ANGTOL � Z
 	 A�   �����PPINFO 6� 5�8�J�\�n���  B�p��� ���������!��E�/�U�{�h��ߧ��� ������%7I�[m��PPLI�CATION ?}���h��LR Ha�ndlingTo�ol � 
V�9.10P/03���
8834�0��
F0�9�51����7�DF1� ��No�ne�FRA�� 6%�_�ACTIVE� � ���  �U_TOMOD�:���ӪCHGAPO�NL� �OUPLED 1^�� * ./@/R/��CUREQ 1	�^�  T\)\,�\,	�/�%� �$�w\"��Ƣ$H�%-"�*H�TTHKY�/��$\�/�/X?"?�/F? d?j?|?�?�?�?�?�? �?�?TOO0OBO`OfO xO�O�O�O�O�O�O�O P__,_>_\_b_t_�_ �_�_�_�_�_�_Loo (o:oXo^opo�o�o�o �o�o�o�oH$6 TZl~���� ��D�� �2�P�V� h�z�������ԏ� @�
��.�L�R�d�v� ��������П�<�� �*�H�N�`�r����� ����̯ޯ8���&� D�J�\�n��������� ȿڿ4����"�@�FπX�j�|ώϠ��#n%T�O�й�DO_CLEAN��1��NM  �� \/ߑߣߵ���b.DSPDRYR8�&�HI�[�@l�3� E�W�i�{���������������MAX@� ����!	')�X��(%"(�PLUG�G �%#�PRC*��BY�]�"����O�����SEGF�K������Y�k߀3EWi{����LAP�#�#��� );M_q�����TOTAL�K�t�#USENU
 + ��/�"n �RGDISPMM�C��;1C��;�@I@�$O�0����#_STRING� 1
�
�kM�S�
~!�_ITEM1�&  n��/�/�/�/�/ �/?"?4?F?X?j?|?��?�?�?�?�?�?�?�I/O SIG�NAL�%Tr�yout Mod�e�%Inp:@S�imulatedލ!OutLL�OVERR� =� 100�"In� cycl@E�!�Prog Abo�rVC�!6DSta�tus�#	Hea�rtbeat�'MH Faul�G�CAler�IO�O __1_C_U_g_y_�_�_ ӄ+і/ �_�_ oo$o6oHoZo lo~o�o�o�o�o�o�o��o 2�_WOR ���+jq�_D��� �����"�4�F� X�j�|�������ď֏�PO�+�A��{ ��1�C�U�g�y����� ����ӟ���	��-��?�Q�c�u���	�DEV���%���ٯ��� �!�3�E�W�i�{��� ����ÿտ�����>/�PALT�]V� �0�~ϐϢϴ����� ����� �2�D�V�h��zߌߞ߰���D�GRI.��+��n���"�4� F�X�j�|������ ��������0�B�T�f����R�]���x� �������� 2D Vhz��������
��PREG Z�C��j|�� �����//0/ B/T/f/x/�/�/�/M��$ARG_jpD ?	����!��  �	$F	[�8]7�G&9� S�BN_CONFIQG@�+DACB>1�CII_SAVE  Dc1Z2� �TCELLSET�UP �*%  OME_IOM�L%MOV_H8�0�?�?REP��O��&UTOBACK�1�)`1F�RA:\0 XO0}0'`�@0>[F � lK_0� 18/�02/09 11�:06:040�'80�O�O_�OLL��'_N_`_r_�_�_�_0�<_�_�_�_oo 0o�_Tofoxo�o�o�o �oKo�o�o,> �obt���������  GA_*C_�\ATBCKCTL.TM����1��C�U�KINIY��0V5$CMESSAGr0|�}1� ��ODE_D�0u6V5�f1��O����$CPA�US�!��+ ?,,		�'0�% �,��L�6�X�Z�l� ����ʟ��Ɵ ��$��� �Z������TSK  �[Oa��'@UPDT��z�d�ˠˆXWZD_�ENBz�R:ԦST�Ay��!˥�!XIS~D0UNT 2�%�c1|0� 	����o��M����ݬ�'�� �C06�{3g��R���v��� ��� ��a3}I}@ʡ�ڿ��׿�.�MET��2��~3� P5�?�UY�?�??B;��50�>�RL�<o��6�D��<�0�<���r��;i�8;����SCRDC�FG 1�%N=A �z5z2�� ������	��-�TO0Qv9��}ߏߡ߳��� ��>���b��1�C�U��g�y�����'*AGR`���ߏ���pNA�0��+	*D��_E�Dx�1��� 
� �%-�pED�T-���:6�Z���Π~E �+B)�0'2�_�6"���  ����2���;��&�t����_����N����3 ��+=�+r����4c�� �=��>P�t��5//�|/�=X/@�/
//�/@/��6�/ k/H?�/=$?�?�/�/~??��7�?7?O[? =�?[O�?�?JO�?��!8�O;��O_��>�O@'_nO�O_�O��9__�O�_�O�>�_�_:_0L_�_p_��CR��O wo�o8MRo�ooo�o�:o���NO_DE�L����GE_UN�USE����IGALLOW 1���   (*SYSTEM*��	$SERV_�GR�{wp��REGƀu$�s�wpNU�M�z�s�}PMU|#p�LAY/���PMPA�Ly��uCYC10�~���=�UL�SU��}����s�LS���BOXOR<İ�sCUR_y��}�PMCNV�v�y�10-�߀T4�DLIߠr��y	*�PROGRAt?PG_MI�/�FA�AL�N�8�A��Bl�w~$FLU?I_RESU����L��l�o�� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2ϕh���LAL_OUT� f{����WD_ABOR�G~�����ITR_RTN�  �T�Py��N�ONSTO����� ��CCG_CONFIG ��L������&�8���E?_RIA_IDp���`�Tq��FCFG ����]�i�_PA��GPw 1s���A�������߾�C�P� �"���C��C �"�("�-�C8"�@�"�H"���CX"�`�"�h"�p"�x䤪"�"�"�"�`������U?����HE�`ӥ���G_mP��1�� 5� s6�$�6�H�Z�l�~����B�HKPAUSf��1��`� -� ����������B (fx^����@���,>�Om��s��WXpCOL_LECT_m���c��uEN�p��Or�NNDE}�����b1�234567890��R�q�����S#
 U�]��Q)0/U/ �l//A/�/�ks/�/�/ �/�/�/&?�/??n? 9?K?]?�?�?�?�?�? �?�?�?FOO#O5O�O�YOkO}O�O�O��q2�� ��IO  ���X��`X_j_|_�_&WTR��S2!
]E� AY
�O�^�"5]�ZHu��_MORR#�� y���Oe 	 Oi goUo�oyo�o�k(b��*Q$6m,Hu?����	�sKPKtKQAR��%PR&�g��Xj|�
I�kр���Q��rZӝ�us �a�PDBT�(���Dcpmi�dbg�T��f�:���N;�p@���d�/  ��N>�ݏ���ܺ���%�����mg�o�:����f^������@u�d1:ܟ��Z�D�EF '@S)��c�buf.�txt�^���_KMC/c)��Sd����.d*��u���ѥ�v�Cz  B*!�`C�ظ�B��0CCI;�p����C;_�Ǻz�`E���D]qeD��J0?M�D�I�>ڐ�
��F��FR���F@��CH��F@��B�q�P�y�b}��g,
\TШk!KP�`KPJ�`��`��T�m����@ Da  �D�  E	� �D�@ ˱2�|� Fp F"�� G=�fF�ߚG'i
�G>��Gg� GK�  H�<=H��&HyMZ���  >�33  `C���n���r�#5YKşbQ�Aq�t=L��<#�e�MQ���Ş|�RSMOFST %/��:HP_T1��D�E -*��X�Qw�KQ;��������?���<�\2��EST)�+/����R.X��զC�4y��z�KPm��{����T�B�R���p���?�KP:d��
��T_)�PROOG �Ʃ�%o��I��.PNUSER�����\�KEY_TOBL  ����h�9��	
�� �!"#$%&'()*+,-./��:;<=>?@A�BC)�GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������#����͓���������������������������������耇����������������������A�LCKg��^�g�STAT����_AUTO_DO�9����IND���btR�����T2*�z�STO�NT{RL�LETE��q
_SCREE�N 6jk�csc�Ub MM�ENU 1/%� <8�7���u� =̓@yPb �������-/ //c/:/L/�/p/�/ �/�/�/�/?�/ ?M? $?6?\?�?l?~?�?�? �?O�?�?OIO O2O OVOhO�O�O�O�O�O �O�O3_
__i_@_R_ x_�_�_�_�_�_�_o �_o,oeo<oNo�oro �o�o�o�o�o�o O&8�\n�����ƙ�_MA�NUALf�DB;CO RIG����&�_ERRL%�	0��X�Eߖ������ C�NUMLI�2�M�����DB�PXWORK 11�����,�>�P�|b�v�DBTB_|G 2r�ѣ��ؤ�	�DB_AWA�YK�X�GCP r��=<ж�_AL2�����G�Ye ���<��_e� 13� , 
	�G���5�r��|�_M I��Ĝ@||���ONTIM���������
�v��MOTNEN���m��RECOR�D 19�� �<z���G�O�B�0� ��Œn�������;��� ӿB���f��-�?�ֿ �u�俙�Ͻ����� �ώ�߆�;ߪ�_�q� �ߕ�߹�(���L�� �%�7��[������ �������H���l�� ��E�W�i�{����� ��2�������A ,:w�����. ��d�=Oa �p��*�� /��9/�]/��/ �/�/�/R/�/J/�/n/�#?5?G?Y?�/��TO�LERENCÔB���ѐL��C�C�SS_CNSTC�Y 2:�����\?
���?�?�?�?O O,O>OTObOtO�O�O �O�O�O�O�O__�4�DEVICE 2;�; ��i_h_ �_�_�_�_�_�_�_o�o{��3HNDGDg <�;7�Cz7n_LS 2=P]/o �o�o�o�o�o�o1o��2PARAM �>#��u\�4SL?AVE ?Pm<g_CFG @9�sdMC:\��0L%04d.CSV
�c�	��"�A �sCH�pba�b�~�-�vW�v��J�Z�H�G���JCP�z�o_
������~tRC_OUT �AP]��_SG�N B��&j���27-F�EB-18 10�:38�p�0=9�1:06�pyV LIX�9��5�~6���+��i��Þ�����I�|uVERSIO�N ��V�4.1.0��EF�LOGIC 1C^�; 	r���ԙ�䝶�PROG�_ENB��Xf�U�LS�� Wf��_�ACCLIM����ss�C�WRSTJN��٥�����MO���ur��I?NIT D�:�v� ��OPT`p� ?	����
 ?	R575s74�6��7��5���1�2��r�B�|��ѤTO  ݭ�L�����V��DEX�p�d{�����PA�TH {�A�\�����s;HCP�_CLNTID y?��qs ���3N�}1IAG_G�RP 2I�y ��� 	 �@K�@G��?���?l��>���dʘ��1���d�����0����?ϧb�?� �i��^?�Vm?S���d�f403� 6789012�345>ғ���� ���s��@n���@i�#@d��/@_�w@Z~��@U/@O��@I��@D(��d�\О�@��tpX�p�ѓ0A�0�0�pB4d�]Pd�ݨꞁ
[�1��-�@)hs@$���@ bN@���@e���@?�D@+������߸Խ��н���R���@N@I��@D�@>�y@9��@4���.v�@(��@"�\�%�7�I�[����L�@Gl��@BJ@<z��@6e�0�`@*�y�$��@�������������=q@q���F@|�@3�3@�R@-�?���?��`?�++�=�O��a�s�����-�@&�@��}��!?�?� ŷ������� ���׋����� ��C!Sy _����	/� /Ţ��p��ш���, ���t!Y��?��?�z�!��o5AF�!4�� ��L4R�!޳�@�p��"�Q���"-� � Q�@��U ��Ah��=H��9=Ƨ�=�^�5=�0��>����=�,v'?�,7� ����C��<(�UC�c 4�¤�k?��d�A@��?��3/�?;- �?�?�?��d4�?)O�?�9O_OAO�O�O?)>���y�B�R=�?��=��z�A��o��G��OG���@�u�uWW�.T@�p�ғ6�̷uB����X B�B�?�B%��͟�$�_p^'Q��U���Q�Q�L�\c���Ѩ*���� B�@B��B��A��@��_c�0o��<~�5o^opo@?�o�oo�ot[�o��bd�C������CgxC޼з����?H�o4�oXC|�g�e�DICT_�CONFIG �J����/��eg��u�STBF/_TTSp�
��sЋ�O�F����MA�Uj���MSW_kCF�pK��  ��~ڊOCVIEW"�3Lb�����Lo�� Ə؏����S���7� I�[�m���� ���ǟ ٟ������3�E�W� i�{�����.�ïկ� ������A�S�e�w� ����*���ѿ���� �+Ϻ�O�a�sυϗ� ��8���������'ߖs�RC[�M�/�! ��5�_ߔ߃߸ߧ������ ��SBL_FAULT NR�|w��GPMSK��-��pTDIAG �O�y�Q'���'�UD1: �67890123�45���r~��w5�P ���������� �2� D�V�h�z���������@������z�5ِ2
��|.�vTRECPc�u�
��u��6�� ����/A Sew��������
/x�UMP_OPTION��&�3!TR[��*��T%PME�G/Y_�TEMP  ï��3B�P� ��Q�$UNI@���!�O�YN_BRK �P��R�EDITCOR9!?!�/�"_K �ENT 1QR��  ,&ST?YLE1 -!/{m&PROG_:?�w?&-BCKEDTh?z?���?�r��?�?�?O�?'O NO5OrOYO�O�O�O�O �O�O_�O&__J_1_ C_�_g_�_�_�_�_�_ �_�_"o4ooXo?o|o��o�pEMGDI_STA�%�q�!�%�NC�c1Rb� ����o�o".
".d 	/L^p���� ��� ��$�6�H� Z�l�~�������Əa% ݏ���!�9q!�G� Y�k�}�������şן �����1�C�U�g� y�������)�֏�� ��0�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ��ί�������(�2� D�V�h�zߌߞ߰��� ������
��.�@�R� d�v�����ϴ��� ��� ��<�N�`�r� �������������� &8J\n�� ���������*� 4FXj|��� ����//0/B/ T/f/x/�/�/���/ �/�/?",?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�/�O�O�O _? $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�O�o �o�o�o_.@R dv������ ���*�<�N�`�r� �����o��̏ޏ��
 &�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφ� ����������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ���������� �2� D�V�h�z��������� ������
.@R dv������ ���*<N`r �������/ /&/8/J/\/n/�/� ��/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�/�/�O�O�O �O�/__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �O�o�o�o�o�O  $6HZl~�� ������ �2� D�V�h�z��o���� ԏ�o��
��.�@�R� d�v���������П� ����*�<�N�`�r� ��~�����̯���� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�jτ����ϲ� ���������0�B� T�f�xߊߜ߮����� ������,�>�P�b� �ώϘ��������� ��(�:�L�^�p��� ������������  $6HZl��� ������ 2 DVhz���� ���
//./@/R/ d/~l/�/�/�/��/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\Ov/�/�O �O�OlO�/�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo TonO�O�o�o�o�o�O �o�o,>Pb t������� ��(�:�L�^�xo�� �������o܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�p�z�������ʏ �����
��.�@�R� d�v���������п� ����*�<�N�h�Z� �ϖϨ�¯ԯ����� �&�8�J�\�n߀ߒ� �߶����������"� 4�F�`�r�|���� ����������0�B� T�f�x����������� ����,>��j� t�������� (:L^p� ������ // $/6/H/bl/~/�/�/ ��/�/�/�/? ?2? D?V?h?z?�?�?�?�? �?�?�?
OO.O@OZ/ HOvO�O�O�/�O�O�O �O__*_<_N_`_r_ �_�_�_�_�_�_�_o�o&o8oRO �$E�NETMODE �1S�E��  b@b@�]Eo�ka`RROR�_PROG %�nj%\F�o�i�eTA�BLE  nk��O 2DRw�bSE�V_NUM }b?  �xatp��a_AUTO_ENB  �evc�dw_NO�q Tnk��asr  *�*�p��p��p��pp�+�p��	��tFLsTR��vHISps�`Av`�{_ALM �1Unk �]D�|\@+
�����ɏ�ۏ����_ir�p  nk�q�bD�a`�TCP_VER �!nj!�o�$E�XTLOG_RE�QE��y��SI�Z����STK����u���TOL � `ADzM��{A ��_BWD$�`��)�%��b�DI�w V�E)�x�d`A*�STEP;��M�a`g�OP_DO�ޟ_aFDR_GR�P 1Wni/�d �	?�ܯ�`͠n&����c?���$,MT�� ��$ ����ͣ"�3��V�A� z�e�����¿����������@��As�>(��#�~b@
 E��`B @�Kϗh>���ϲϝ������A@f���@�/33@���Ӽ́@��߻�D�V�͠F@ l�`�`�l�\���L�FZ!D��`�D�� BT��@���4��?�  ��Z�6��������5�?Zf5�ES��4���@��`O������a�Y`����+�kFEATUROE X�E%��a�LR Ha�ndlingTo�ol ^�`BE�nglish D�ictionar}ya�4D StS��ard^�`�Analog I/O�����gle Shi�ft��uto S�oftware �Update��m�atic Bac�kup_��gro�und Edit�W�a�Camera���F��Commo�n calib �UI8�D�n�O�M�onitor\�t�r\�Reliab<��`�DHCP9�^��Data Acq�uisk��iag�nos����oc�ument Vi�ewew��ual� Check S�afetyW�d�hancedW�`�-�s  Fr0�b�xt�. DIO g�f�i��\end1 E�rrv�L��xPs�w	r��g  �^�F�CTN Menu� v���TP I�n� fac�c�G��p Mask �Exc- gYHT�� Proxy S�vigh-S;pe1 Ski����k mmunicn��onsVur� � �����conn�ect 2�nc=r� struu�_��KAREL Cmod. Lua~�Run-TiX �Env�� el u+ �s��S/Wa�License� � Book(S�ystem)^�M�ACROs,M/�Offse��T%H0k ���Y MRp�l���M����l MechStop+t���T%i����&ax1 �����.od��witch?�#��y.y&4;OptmF?L�#,fi�.�&g�~T%ulti-T�"�_�PCM fu�n��9a� tiz��8�7o��Regi�I rq�6ri��F��;F��Num S�el�%/IV  Ad�jua*NWA��hMt�atuA�O��c�R�DM Robot>r�scove{�Eem� kn��E�BServok !0`�?SNPX b"��;SN� Cli��#^��Librz�C_S�Q �$UPVo. t� �ssag�5d�X� 0��l!��X�/I��U�MILIB�_�RP� Firm��^P��Acc�!�TPsTX���Telnl ��_�Q[�h%�]orq}u��imulau�6�U��B3&+e3v.�U��ri 8o�Unexcep	t1 �@n�eQ��VCS�rlc�(V@��r o*uU[${S6PsSC2e\SUI��?Web Pl�F�~�Q��t3+��ZDT Applj�^�iP� a<Y� �Grid�Apla�y��P��Rr.���X���1"� ��2�00i���sciyi+VBLoad  ��Upl;���gPat)6(�yc��`�@�` �RL��V �y MI Dev$  (QM"�6���7sswo���/�64MB DRA9M���FRO��-�gell��B�sh̑�؟�ce;���pa\
!�sty��sAB��t�^0.���@kX���6� 2�a��port?�@ R��q$T1p�	[� ��d�No m�@{�c��d�OL[�Supx��}1HOPT ��,�Z�S� cro��L�CUUL��NF���uWestUS[�e�'texqdUp�Ư_PP� %OToeu(0P+�s{rt|�C�stdpn�k�s� SWIMES7T fv�F0]�b��W��i�{Ϩϟϱ� ���������7�A� n�e�wߤߛ߭����� �����3�=�j�a� s����������� ��/�9�f�]�o��� ������������ +5bYk��� ����'1 ^Ug����� � /�	/#/-/Z/Q/ c/�/�/�/�/�/�/�/ �/??)?V?M?_?�? �?�?�?�?�?�?�?O O%OROIO[O�OO�O �O�O�O�O�O�O_!_ N_E_W_�_{_�_�_�_ �_�_�_�_ooJoAo So�owo�o�o�o�o�o �o�oF=O| s������� ��B�9�K�x�o��� �������ۏ��� >�5�G�t�k�}����� ����ן���:�1� C�p�g�y�������ܯ ӯ���	�6�-�?�l� c�u�������ؿϿ� ���2�)�;�h�_�q� �ϕϧ���������� .�%�7�d�[�mߚߑ� ������������*�!� 3�`�W�i������ ��������&��/�\� S�e������������� ����"+XOa �������� 'TK]�� ������// #/P/G/Y/�/}/�/�/ �/�/�/�/???L? C?U?�?y?�?�?�?�? �?�?O	OOHO?OQO ~OuO�O�O�O�O�O�O ___D_;_M_z_q_ �_�_�_�_�_�_
oo o@o7oIovomoo�o �o�o�o�o�o< 3Eri{��� �����8�/�A� n�e�w�������Ǐя �����4�+�=�j�a� s�������ß͟��� �0�'�9�f�]�o��� ������ɯ�����,� #�5�b�Y�k������� ��ſ����(��1� ^�U�gϔϋϝϷ��� ������$��-�Z�Q� cߐ߇ߙ߽߳����� �� ��)�V�M�_�� ������������ �%�R�I�[������ ����������! NEW�{��� ���JA S�w����� �///F/=/O/|/ s/�/�/�/�/�/�/? ??B?9?K?x?o?�? �?�?�?�?�?O�?O >O5OGOtOkO}O�O�O �O�O�O_�O_:_1_ C_p_g_y_�_�_�_�_��_ o�_	o6o-a � H551�+cQa2VfR782�Wg50WeJ614�WeATUP{f54�5{h6WeVCAM�WeCUIF{g28n�fNREcf52�fwR63bgSCHWe�DOCV�fCSU�cf869{g0�fE�IOC�g4nfR6=9�fESET�g�g{J7�gMASKWe�PRXY�h7WfOCO_x3�hnfgpzh�yh53"vH�xLC�H�vOPLG�g0^�vMHCR�vS�wMAT�fMCS�h�0jw55�fMDS�W[��wOP�wMP�R�v�`�v+pzfPCM�g5��gp�f���[51�g51҈0�f�PRS^w69�vF{RD�fRMCNWf{93zfSNBA�g^�wSHLB3�MU�t�`N�2zfHTC�f�TMILch"vTP�A:vTPTX��E�L&��"w8mgJ9�5�fTUT�vUE�C�vUFR�fVCuC
�O�VIP���CSC��pIWeW�EB�fHTT�fR�6�hؘCG]�IG�E�IPGS��RCv��DG�wH75�f�R7QwRЈR66ڲx2�vR6UgR5�5�4Vf�`VfD0u6�fF(�CLI����gCMS:vW��fS[TY.�TO^�7!w��`�fORS�R6u8zfM �NOM:v�OLA�OPI��SWENDcfL�S���ETS��+p��CPv�g78VfFVR:v�IPN��Gene Wd2h]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'��9�  H�551;�U�2Z�R�782[�50[�J�614[�ATUP���545��6[�V�CAM[�CUIFv��28��NREk�52��R63j�S{CH[�DOCV;�wCSUk�869��0��EIOC�4�z�R69��ESE�T����J7��MA{SK[�PRXY��]7[�OCO��3��z������53j�H�HLCH��OPL�G��0*
MHCR���S�MAT
�MkCS��0��55���MDSWOPMPR
'�

w�.��PCM��5i��ؚ� Z51��51��0��PRS��6�9

FRD��RM�CN[�93��SN�BA�ISHLB�+*MY+'��2��H{TC��TMILk��j�TPA��TPT�X�*EL*� j�8�y�J95��TUT�
UEC��UFR���VCCJ<O�
V;IP�*CSC�*X��I[�WEB��HT�T��R6�<CG��;IG�;IPGS��:RC�*DGH[75��R7��R��R66*2*
R6.Y�R55zL4Z��Z�D06��F�LCsLIJ��CMS���P��STYz;TO�;7i����ORS��
R68��M�N�OM��OL�OP�I
JSENDk�L:Y;Sh\ETS
Jw�+CP
�78Z�F�VR��IPN�*Gene[�:�aoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%��7�C�STD~>�LANG_� Z�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx��� ����//,/>/�P/b/t/�/�/�*RB=T^�OPTN�/�/��/�/?DPN ]�-???Q?c?u?�?�? �?�?�?�?�?OO)O~;Oted _� 6�eOwO�O�O�O�O�O �O�O__+_=_O_a_ s_�_�_�_�_�_�_�_ oo'o9oKo]ooo�o �o�o�o�o�o�o�o #5GYk}�� �������1� C�U�g�y��������� ӏ���	��-�?�Q� c�u���������ϟ� ���)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�9�K�]�o��� �������������� #5GYk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_  ��_�_�_�_o� o2m999e�$�FEAT_ADD ?	���fa�n`  	 6hwo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/�5/G/Y/YdDEMO� Xfi   6h�-�/�/�/�/ �/???A?8?J?d? n?�?�?�?�?�?�?O �?O=O4OFO`OjO�O �O�O�O�O�O_�O_ 9_0_B_\_f_�_�_�_ �_�_�_�_�_o5o,o >oXobo�o�o�o�o�o �o�o�o1(:T ^������� � �-�$�6�P�Z��� ~�������Ə���� )� �2�L�V���z��� ��������%�� .�H�R��v������� ������!��*�D� N�{�r���������� ޿���&�@�J�w� nπϭϤ϶������� ��"�<�F�s�j�|� �ߠ߲��������� �8�B�o�f�x��� �����������4� >�k�b�t��������� ����0:g ^p������ 	 ,6cZl ������/� /(/2/_/V/h/�/�/ �/�/�/�/?�/
?$? .?[?R?d?�?�?�?�? �?�?�?�?O O*OWO NO`O�O�O�O�O�O�O �O�O__&_S_J_\_ �_�_�_�_�_�_�_�_ �_o"oOoFoXo�o|o �o�o�o�o�o�o�o KBT�x�� �������G� >�P�}�t��������� ������C�:�L� y�p����������ܟ ���?�6�H�u�l� ~��������د�� �;�2�D�q�h�z��� ����ݿԿ� �
�7� .�@�m�d�vϣϚϬ� ���������3�*�<� i�`�rߟߖߨ����� �����/�&�8�e�\� n������������ ��+�"�4�a�X�j��� ��������������' 0]Tf��� �����#, YPb����� ���//(/U/L/ ^/�/�/�/�/�/�/�/ �/??$?Q?H?Z?�? ~?�?�?�?�?�?�?O O OMODOVO�OzO�O �O�O�O�O�O_
__ I_@_R__v_�_�_�_ �_�_�_oooEo<o No{oro�o�o�o�o�o �oA8Jw n������� ��=�4�F�s�j�|� ������̏֏���� 9�0�B�o�f�x����� ��ȟҟ�����5�,� >�k�b�t�������į ί����1�(�:�g� ^�p���������ʿ�� � �-�$�6�c�Z�l� �ϐϢϼ��������� )� �2�_�V�hߕߌ� �߸���������%�� .�[�R�d����� ��������!��*�W� N�`������������� ����&SJ\ �������� "OFX�| ������// /K/B/T/�/x/�/�/ �/�/�/�/???G? >?P?}?t?�?�?�?�? �?�?OOOCO:OLO yOpO�O�O�O�O�O�O 	_ __?_6_H_u_l_ ~_�_�_�_�_�_o�_ o;o2oDoqohozo�o �o�o�o�o�o
7 .@mdv��� �����3�*�<� i�`�r�����Ï��̏ �����/�&�8�e�\� n���������ȟ��쟀��+�"�4�a�X���  {������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^ p�������  $6HZl~ �������/  /2/D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�o 0BTfx��� ������,�>� P�b�t���������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l�~� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� ��������*�<�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^/|p/�)  �( �!�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�o�o 0BTfx� �������� ,�>�P�b�t������� ��Ώ�����(�:� L�^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ������¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���������*� <�N�`�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j� |��������������� 0BTfx� ������ ,>Pbt��� ����//(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�?�? �?O O2ODOVOhOzO �O�O�O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo*o <oNo`oro�o�o�o�o �o�o�o&8J \n������ ���"�4�F�X�j� |�������ď֏��� ��0�B�T�f�x��� ������ҟ����� ,�>�P�b�t������� ��ί����(�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ������� ��� �2�D�V�h�z� �ߞ߰���������
� �.�@�R�d�v��� �����������*� <�N�`�r��������� ������&8J \n������ ��"4FXj |������� //0/B/T/f/x/�!� (�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x�����$FEAT_�DEMOIN  ������������INDEX��������ILECO�MP Y����������SETUP2 �Z���� � N %��_AP2BCK 1[�?  �)��Y�"h�%O������z� ����N��r�ϖ�� =�̿a��ϗ�&ϻ� J����π�ߤ�9�K� ��o��ϓ�"ߠ���X� ��|��#��G���k� }���0�����f��� �����,�U���y�� ����>���b���	�� -��Qc���� :��p�); �_���$�H ��~/�7/�D/ m/��/ /�/�/V/�/ z/?!?�/E?�/i?{? 
?�?.?�?R?�?�?�? O�?AOSO�?wOO�O �O<O�O`O�O_�O+_��OO_�O\_�_��3�P�7� 2L�*.cVR�_�_DP*�_��_ASo)oU�PPC�1oZoDPFR6:DEo�no�o9kTΠ �o�ooe�o
|���o0V*.F�_aCQ	qcO�|�A{STM �r��nt`���DPiPe�ndant Pa'nel�A{H�i���wW�����BzGIFŏ��uۏ����?�BzJPGI�s��u_�0�.�ß:jJS͟���DP��䟡�%
J�avaScript"�M�CS�z��v�g�$� %Cas�cading S�tyle She�ets��P
AR�GNAME.DTկ8\�p\鯧�	���*�֯�DISP* ���pm���<������Z�	PANE3L1���%�p�1�$�6��2&ό�� z�7�I����3���@��ϻ���b��4.߀��ǂ�?�Q����T�PEINS.XML�߉�:\�����Custom T?oolbarB�a��PASSWORD���6^FRS:\���D� %Pas�sword Config��_��� �E�k_i������.� ��R���������A ����w�*�� `��+�O� s��8�\n /�'/� /]/��/ /�/�/F/�/j/�/? �/5?�/Y?�/�/�?? �?B?�?�?x?O�?1O CO�?gO�?�O�O,O�O PO�OtO�O_�O?_�O 8_u__�_(_�_�_^_ �_�_o)o�_Mo�_qo  oo�o6o�oZo�o �o%�oI[�o ��D�h��� 3��W��P������ @�Տ�v����/�A� Џe�􏉟�*���N� �r�ܟ���=�̟a� s����&���ͯ\�� �������K�گo��� h���4�ɿX������ #ϲ�G�Y��}�ϡ� 0�B���f��ϊ���1� ��U���yߋ�߯�>� ����t�	��-���� c��߇����L��� p�����;���_�q��O��$FILE_�DGBCK 1[���X���� < �)�
SUMMARY�.DGu�!�MD�:����-�Di�ag Summa�ry����
CONSLOG������-�m��Conso?le logn��	TPACCNc��%����TP� Account�in���FR6�:IPKDMP.'ZIP!%�
9r���	Except�ionv��*.�DT��-�FR�:\���FR� DT File�s�&��MEMCHECK�J��}/��Memory� Data~/M���`�)	FTP�`�/d/�/�'�m�ment TBD�?M�L >))�ETHERNET��/�<!E?�?��E�thernet ~� figura�����!DCSVRF��/�/�/O�!%��0 verify� all
OO�M{,�5DIFF�?p�?�?�O� %!Hdiff�OBG<!�0CHG01�OjO|O`_A�O9_DB*��I2_�O _�_�O6_H_��B3�_r_�_o ��_@o�VVTR�NDIAG.LS�Eo�_o�o�!]a �Ope�3 Log� nostic�M�T4�)V7DEVabDA�zox�o!AVis�a?Device�o�kIMGabh�o�z�S9tImagEn�kUP�`ES�o~~FRS:\�����Update?s List*�����pFLEXEV�EN{?����A�p� UIF Ev�1�`��  +�l�)
PSRBW�LD.CMُ!����,�� PS_R?OBOWEL#?��}��HADOW����������#Sha�dow Chan�g/�&�L�s�RCMERR�������7��#��CFG �Error?pta�ilڟ S�|;"��SGLIB/���(����!�� S�t�0�ad�u��)��ZD�/���;�n�'ZD�`adݯzj�r�NOTI�?��,����%Not�ific�2j�ㆀAG��'�<�K�I� r����%Ϻ���[��� ��&ߵ�J���n߀� ߤ�3���W����ߍ� "��F�X���|��� ��A���e������0� ��T���a������=� ����s���,>�� b����'�K� o��:�^p ��#��Y�} /$/�H/�l/�y/ �/1/�/U/�/�/�/ ? �/D?V?�/z?	?�?�? ??�?c?�?�?O.O�? RO�?vO�OO�O;O�O �OqO_�O*_<_�O`_ �O�__�_�_I_�_m_ oo�_8o�_\ono�_ �o!o�o�oWo�o{o �oF�oj�o�� /�S����� B�T��x����+��� ҏa������,���P� ߏt������9�Ο�� o����(���5�^�� �������G�ܯk� � ���6�ůZ�l����� ���C����y�ϝ� 2�D�ӿh����Ϟ�-� ��Q����χ�߫�@� ��M�v�ߚ�)߾��� _��߃��*��N����r���$FILE�_FRSPRT � ��h�������MDONLY 1[��~_� 
 �� ��7��[��D��h� �����-���Q����� ����@R��v �)��_�� *�N�r�� 7��m/�&/� 3/\/��//�/�/E/ �/i/�/?�/4?�/X? j?�/�??�?A?�?�?~��VISBCK��|����*.VD�?|9O�0FR:\@�ION\DATA�\$O�2�0Vi�sion VD fileeOs?�O�O �?�O�?_�O_=_�O a_�O�_�_&_�_J_�_ n_�_o�_9oKoooo �_�o"o�o�oXo�o|o #�oG�ok�o �0������ �0�U��y������ >�ӏb�������-����LUI_CONF�IG \��|A8� $ ���{�叟����şן���w�|x�!�3� E�W�i�y�������� ү�{����,�>�P� b�����������ο� w���(�:�L�^��� �ϔϦϸ�����s� � �$�6�H�Z���~ߐ� �ߴ�����o���� � 2�D�V���z���� ����k���
��.�@� ��Q�v���������U� ����*<��` r����Q�� &8�\n� ���M���/ "/4/�X/j/|/�/�/ �/I/�/�/�/??0? �/T?f?x?�?�?3?�? �?�?�?OO�?>OPO bOtO�O�O/O�O�O�O �O__�O:_L_^_p_ �_�_+_�_�_�_�_ o o�_6oHoZolo~o�o 'o�o�o�o�o�o�o 2DVhz�#� �����	�.�@� R�d�v��������Џ �􏋏�*�<�N�`� r�	�������̟ޟ� ���&�8�J�\�n�� ������ȯگ쯃�� "�4�F�X�j����������Ŀֿ�x��x���  �$FLU�I_DATA �]���-���RESU_LT 2^-�V�� �T�/�wizard/g�uided/st�eps/Expertύϟϱ����π������/�A�O���Continu�e with Gj�anceOߊߜ� ������������,�,>�P� �-�-�>o�0 ���o��/�.����a�ps R��������"�4�F� X�j�|�����_Є��� ������!3EW i{�������:����ripx��� );M_q��� ������/%/7/ I/[/m//�/�/�/�/ �/�/�/��?������s�TimeUS/DST?�?�? �?�?�?�?�?OO/O�AOX�Disablx�vO�O�O�O�O�O��O�O__*_<_N^
�{�7?)?;?M?_?q224x?�_�_o o%o7oIo[omoo�o PObO�o�o�o�o! 3EWi{��^_�p_�_�_�_�_zon u0�5�G�Y�k�}��������ŏ׏�X�E�ST Eap�rn? Stande�� ,�>�P�b�t�������`��Ο���a� �{�������`�r�acces������ ��̯ޯ���&�8��S�c�nect �to NetworkG�~�������ƿ ؿ���� �2�D��a��!���E��!Y��o0IntroductionJ����� ��'�9�K�]�o߁� ��/����������� #�5�G�Y�k�}����?qϻ��  ���s/Safety��-�?�Q�c�u��� ������������ );M_q��� �����r����8����e�Reg��~ �������/� /2/��Europ�om//�/�/�/�/��/�/�/?!?3?E?zc�?AS�EUF?�?�?�?O!O�3OEOWOiO{O�O��C|	�X"an Ce��al�O�O�O�O__ *_<_N_`_r_�_�_U6��?u?�?�?�?� "�'o9oKo]ooo�o�o �o�o�o�o���o# 5GYk}��� ��� �_�_�_�_|oa/curr�@ ���������͏ߏ����'�9�T�14-�FEB-18 05:03 PM?� v���������П��� ��*�<��R�W+���/�A�S�e�YearB�֯�����0��B�T�f�x����f2018����ο�� ��(�:�L�^�pς��� 
U�o�  ��o��ϓ���c�Month��+�=�O�a� s߅ߗߩ߻������e2����1�C�U� g�y���������� �϶�a3��������g�Day��}������� ��������1�g14;bt�� �����(:����y;�M�c�Houį��� //+/=/O/a/s/�/��5�/�/�/�/�/�/ ?!?3?E?W?i?{?�?L
�k�?���inute�?(O:O LO^OpO�O�O�O�O�O�O��3�O	__-_?_ Q_c_u_�_�_�_�_�_�_�?
��?!o�?�?c�AMc�xo�o�o�o �o�o�o�o,C	 go\n����������"�4�L�L���c�o+o=oOl�NetMethod:�̏ޏ����&��8�J�\�n�����N�ot configure����ϟ� ���)�;�M�_�q������TV�h�z��� ����)�;�M�_��q���������˿ݿ  ���&�8�J�\�n� �ϒϤ϶������U��ͯ��ï%��L�^� p߂ߔߦ߸�������  ��$��H�Z�l�~� �������������  �2�����w�9ߞ� ����������
. @Rdv5��� ���*<N `r�C��g���� �//&/8/J/\/n/ �/�/�/�/�/�/��/ ?"?4?F?X?j?|?�? �?�?�?�?��?�O �BOTOfOxO�O�O�O �O�O�O�O__,_�/ P_b_t_�_�_�_�_�_ �_�_oo(o�?IoO mo/O1o�o�o�o�o�o  $6HZl~ =_�������  �2�D�V�h�z�9o�� ]o��я���
��.� @�R�d�v��������� П�����*�<�N� `�r���������̯�� Տ����#��J�\�n� ��������ȿڿ��� �"��F�X�j�|ώ� �ϲ����������� ݯ'��K�u�7��߮� ����������,�>� P�b�t�3Ϙ����� ������(�:�L�^� p�/�A�S�e�������  $6HZl~ ��������  2DVhz�� ���������/�� @/R/d/v/�/�/�/�/ �/�/�/??�<?N? `?r?�?�?�?�?�?�? �?OO&O��	/kO -/�O�O�O�O�O�O�O _"_4_F_X_j_)?{_ �_�_�_�_�_�_oo 0oBoTofoxo7O�o[O �oO�o�o,> Pbt����� �o���(�:�L�^� p���������ʏ�o� �o��o6�H�Z�l�~� ������Ɵ؟����  ��D�V�h�z����� ��¯ԯ���
��ۏ =���a�#�%������� п�����*�<�N� `�r�1��ϨϺ����� ����&�8�J�\�n� -���Q����߉����� �"�4�F�X�j�|�� ������������ 0�B�T�f�x������� ����ߣ�����> Pbt����� ����:L^ p�������  //����?/i/+ �/�/�/�/�/�/�/?  ?2?D?V?h?'�?�? �?�?�?�?�?
OO.O @OROdO#/5/G/Y/�O }/�O�O__*_<_N_ `_r_�_�_�_�_y?�_ �_oo&o8oJo\ono �o�o�o�o�o�O�O�O �O4FXj|� ��������_ 0�B�T�f�x������� ��ҏ������o�o �o_�!��������Ο �����(�:�L�^� �o�������ʯܯ�  ��$�6�H�Z�l�+� ��O���s�ؿ����  �2�D�V�h�zόϞ� ����ӿ����
��.� @�R�d�v߈ߚ߬߾� }��ߡ��ſ*�<�N� `�r��������� ������8�J�\�n� ���������������� ��1��U�� ������ 0BTf%���� ����//,/>/ P/b/!�/E�/�/} �/�/??(?:?L?^? p?�?�?�?�?w�?�?  OO$O6OHOZOlO~O �O�O�Os/�/�/�O_ �/2_D_V_h_z_�_�_ �_�_�_�_�_
o�?.o @oRodovo�o�o�o�o �o�o�o�O_�O3 ]_������ ���&�8�J�\�o ��������ȏڏ��� �"�4�F�X�); M��q֟����� 0�B�T�f�x������� m�ү�����,�>� P�b�t���������{� �����ß(�:�L�^� pςϔϦϸ�������  ߿�$�6�H�Z�l�~� �ߢߴ���������� Ϳ߿�S��z��� ����������
��.� @�R��c��������� ������*<N `�C�g��� �&8J\n �������� /"/4/F/X/j/|/�/ �/�/q�/��/�? 0?B?T?f?x?�?�?�? �?�?�?�?O�,O>O PObOtO�O�O�O�O�O �O�O_�/%_�/I_? _�_�_�_�_�_�_�_  oo$o6oHoZoO~o �o�o�o�o�o�o�o  2DV_w9_� �qo���
��.� @�R�d�v�������ko Џ����*�<�N� `�r�������g�� ՟���&�8�J�\�n� ��������ȯگ��� ��"�4�F�X�j�|��� ����Ŀֿ������ ݟ'�Q��xϊϜϮ� ����������,�>� P��t߆ߘߪ߼��� ������(�:�L�� �/�Aϣ�e�������  ��$�6�H�Z�l�~� ����a���������  2DVhz�� �o������. @Rdv���� �����/*/</N/ `/r/�/�/�/�/�/�/ �/?���G?	n? �?�?�?�?�?�?�?�? O"O4OFO/WO|O�O �O�O�O�O�O�O__ 0_B_T_?u_7?�_[? �_�_�_�_oo,o>o Poboto�o�o�o�_�o �o�o(:L^ p���e_��_� �_�$�6�H�Z�l�~� ������Ə؏����o  �2�D�V�h�z����� ��ԟ������ =���v��������� Я�����*�<�N� �r���������̿޿ ���&�8�J�	�k� -��ϡ�e��������� �"�4�F�X�j�|ߎ� ��_����������� 0�B�T�f�x���[� ���������,�>� P�b�t����������� ������(:L^ p������� ������E�l~ �������/  /2/D/h/z/�/�/ �/�/�/�/�/
??.? @?�#5�?Y�? �?�?�?OO*O<ONO `OrO�O�OU/�O�O�O �O__&_8_J_\_n_ �_�_�_c?u?�?�_�? o"o4oFoXojo|o�o �o�o�o�o�o�O 0BTfx��� �����_�_�_;� �_b�t���������Ώ �����(�:��oK� p���������ʟܟ�  ��$�6�H��i�+� ��O���Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚ�Y��� }��ϡ���*�<�N� `�r߄ߖߨߺ����� �߯��&�8�J�\�n� ������������ ���1�����j�|��� ������������ 0B�fx��� ����,> ��_!���Y�� ��//(/:/L/^/ p/�/�/S�/�/�/�/  ??$?6?H?Z?l?~? �?O�s�?�?�O  O2ODOVOhOzO�O�O �O�O�O�O�/
__._ @_R_d_v_�_�_�_�_ �_�_�?�?�?o9o�? `oro�o�o�o�o�o�o �o&8�O\n �������� �"�4��_oo)o�� Mo��ď֏����� 0�B�T�f�x���I�� ��ҟ�����,�>� P�b�t�����W�i�{� ݯ����(�:�L�^� p���������ʿܿ��  ��$�6�H�Z�l�~� �Ϣϴ������ϩ��� ͯ/��V�h�zߌߞ� ����������
��.� �?�d�v����� ��������*�<��� ]�߁�Cߨ������� ��&8J\n ��������� "4FXj|� M��q�����// 0/B/T/f/x/�/�/�/ �/�/�/�??,?>? P?b?t?�?�?�?�?�? �?�O�%O��?^O pO�O�O�O�O�O�O�O  __$_6_�/Z_l_~_ �_�_�_�_�_�_�_o  o2o�?SoOwo�oM_ �o�o�o�o�o
. @Rdv�G_�� �����*�<�N� `�r���Co�ogo��ۏ �o��&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯��ߏ��� -��T�f�x������� ��ҿ�����,�� P�b�tφϘϪϼ��� ������(����� ��A��߸�������  ��$�6�H�Z�l�~� =Ϣ�����������  �2�D�V�h�z���K� ]�o�������
. @Rdv���� ����*<N `r������ ������#/��J/\/n/ �/�/�/�/�/�/�/�/ ?"?�3?X?j?|?�? �?�?�?�?�?�?OO 0O�QO/uO7/�O�O �O�O�O�O__,_>_ P_b_t_�_�O�_�_�_ �_�_oo(o:oLo^o po�oAO�oeO�o�O�o  $6HZl~ ������_��  �2�D�V�h�z����� ��ԏ�o���o��o ݏR�d�v��������� П�����*��N� `�r���������̯ޯ ���&��G�	�k� }�A�����ȿڿ��� �"�4�F�X�j�|�;� �ϲ����������� 0�B�T�f�x�7���[� ���ߑ�����,�>� P�b�t������� ������(�:�L�^� p��������������� ����!��HZl~ �������  ��DVhz�� �����
//�� ����s/5�/�/�/ �/�/�/??*?<?N? `?r?1�?�?�?�?�? �?OO&O8OJO\OnO �O?/Q/c/�O�/�O�O _"_4_F_X_j_|_�_ �_�_�_�?�_�_oo 0oBoTofoxo�o�o�o �o�o�O�O�O�O> Pbt����� �����_'�L�^� p���������ʏ܏�  ��$��oE�i�+ ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v�5���Y��� }������*�<�N� `�rτϖϨϺ��ϋ� ����&�8�J�\�n� �ߒߤ߶��߇��߫� �Ͽ��F�X�j�|�� ������������� ��B�T�f�x������� ����������; ��_q5����� ��(:L^ p/�������  //$/6/H/Z/l/+ uO�/�/��/�/?  ?2?D?V?h?z?�?�? �?�?��?�?
OO.O @OROdOvO�O�O�O�O }/�/�/�O_�/<_N_ `_r_�_�_�_�_�_�_ �_oo�?8oJo\ono �o�o�o�o�o�o�o�o �O�O�O_g)_� �������� 0�B�T�f�%o������ ��ҏ�����,�>� P�b�t�3EW��{ �����(�:�L�^� p���������w�ܯ�  ��$�6�H�Z�l�~� ������ƿ������� ͟2�D�V�h�zόϞ� ����������
�ɯ� @�R�d�v߈ߚ߬߾� ��������׿9��� ]�τ�������� ����&�8�J�\�n� �������������� "4FXj)� M�q���� 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/{ �/�?��/:?L?^? p?�?�?�?�?�?�?�?  OO�6OHOZOlO~O �O�O�O�O�O�O�O_ �//_�/S_e_)O�_�_ �_�_�_�_�_
oo.o @oRodo#O�o�o�o�o �o�o�o*<N `_i_C_��y_� ���&�8�J�\�n� ��������uoڏ��� �"�4�F�X�j�|��� ����q��ߟ	�� 0�B�T�f�x������� ��ү����Ǐ,�>� P�b�t���������ο ���ß՟���[� ��ϔϦϸ�������  ��$�6�H�Z��~� �ߢߴ����������  �2�D�V�h�'�9�K� ��o�������
��.� @�R�d�v�������k� ������*<N `r����y�� �����&8J\n �������� ��/4/F/X/j/|/�/ �/�/�/�/�/�/?� -?�Q?x?�?�?�? �?�?�?�?OO,O>O PObOs?�O�O�O�O�O �O�O__(_:_L_^_ ?_A?�_e?�_�_�_  oo$o6oHoZolo~o �o�o�osO�o�o�o  2DVhz�� �o_��_��_�.� @�R�d�v��������� Џ����o*�<�N� `�r���������̟ޟ ���#��G�Y�� ��������ȯگ��� �"�4�F�X��|��� ����Ŀֿ����� 0�B�T��]�7��ϫ� m���������,�>� P�b�t߆ߘߪ�i��� ������(�:�L�^� p����eϯω��� ���$�6�H�Z�l�~� ����������������  2DVhz�� ����������� ��O�v���� ���//*/</N/ r/�/�/�/�/�/�/ �/??&?8?J?\? -?�?c�?�?�?�? O"O4OFOXOjO|O�O �O_/�O�O�O�O__ 0_B_T_f_x_�_�_�_ m??�?�_�?o,o>o Poboto�o�o�o�o�o �o�o�O(:L^ p�������  ��_!��_E�ol�~� ������Ə؏����  �2�D�V�g�z����� ��ԟ���
��.� @�R��s�5���Y��� Я�����*�<�N� `�r�������g�̿޿ ���&�8�J�\�n� �ϒϤ�c��χ��ϫ� ��"�4�F�X�j�|ߎ� �߲��������߹�� 0�B�T�f�x���� ������������;� M��t����������� ����(:L� p�������  $6H�Q�+� u�a�����/  /2/D/V/h/z/�/�/ ]�/�/�/�/
??.? @?R?d?v?�?�?Y� }�?�?�O*O<ONO `OrO�O�O�O�O�O�O �O�/_&_8_J_\_n_ �_�_�_�_�_�_�_�?�?�?�?CoC�$F�MR2_GRP �1_Ke�� �C4  �B�P	 Px�o�l�`F@ �e�E���b�a�Z�a��L�FZ!D��`�D�� BT���@����m?ǀ  �\�`6����)r��5�?Zf5�ES9q�m�A�  Qc{BH�Kt�`}q@�33@%��p�s�\�d��}�`@�q��n�
���a<�z�<����=7�<�
�;;�*�<����m8ۧ�9k�'V8��8����7ג	8(���r��o������̏����W_b_CF/G `lkT�b,��>�P�b��NO �lj
F0�� ����RM_CHK?TYP  \aPpt`v`,`^aROM���_MIN��S������pX_`SS�B�aKe �f�U�0��B��TP_DEF�_OW  T|tcW�IRCOM���h��$GENOV_RD_DOؖQn��THRؖ d���d��_ENB�� ���RAVCecb:��� ��eH�3��W��le�v��z� ���OUh`h�ll���hl��e<������|5�SC�  D^��d�׶Ϗ�@�av�B�Ța|iعI���SMTeci	�x`�Z��$HOSTC�s1jli��_��` MCTr��0�V  27�.0��1i�  e`߭߿������ڛ߀�&�8�J�m����	�anonymou�sq��������� /߄`����^�`�M� ��q��������� ��� ��6���~�[m ����8� �� 4V�EWi{�� �����
@R //A/S/e/w/��� ���/*??+?=? O?�s?�?�?�?�?�/ /�?OO'O9OKO�/ �/�/�O�?�O�/�O�O �O_X?5_G_Y_k_}_ �O"_�?�_�_�_�_o TOfOxO�O�_yo�O�o �o�o�o�o,_	- ?Qto�_�_��� ��(o:oLo)�`M� �oq�������nd�ݏ ���6�7�~[�m� �������� �"� ��V�3�E�W�i�{� ����ïկ�
�@�R��/�A�S�e�w����E�NT 1k�� sP! ���  �����ؿ�п1��� U��a�<ϊϯ�r��� ���Ϻ����?��� u�8ߙ�\߽߀��ߤ� �����;���_�"�� F�|��������� %���1��Z��B��� f��������������Ei,�P
QUICC0�v���1���9��2:(�!ROUTER�fx��!PCJOG���!192�.168.0.1�0��CAMPRYT*//!%1# Q/8&RT�U/g/�/���NAME !~��!ROBOC/��/S_CFG 1�j�� ��Auto-st�artedєFTPܟa1����? )��?�?�?�?�?��O .O@OROu?cO	O�O�O �O�O�O��:?L?^?;_ rO�?R_�_�_�_�_�O �_�_oo%oH_�_[o moo�o�o�o��̟ޟ �4o!h_EWi{ �To����� �/�A�S�e�w����o �o�oя���<�+� =�O��s��������� ޏ`�ڟ��'�9�K� ������ȏʟ����ۯ ����#��G�Y�k� }�����4�ſ׿��� ��f�x���gϞ��� ү�������Ϭ���� -�?�Q�t�u�ߙ߫� ������(�:�L�^�`� 2��q������ ������%�H���[� m����������� � ��4�!h�EWi{ �T�����
 �/ASew?� _ERR l�*���PDUSIZW  ^6 ���>�WRD ?�(5���  guest�//+/=/O/a/�$S�CD_GROUP� 3m(< ,1�"IFT�.$PA�.OMP�. n�._SH�.ED�/w $C�.COM��TTP_AUTH� 1n� <!�iPendan�m'x>#;-Q!KAREL:*x?�?�=KC�?�?�?��0VISION SET� (O�?,V!?O-OWO�3{OiO�O �O�O�O�O_�O�NG4CTRL o��aX
qQF�FF9E3_���FRS:DEFA�ULT�\FA�NUC Web ?Server�ZtQ �J1�$/\�_
oo�.o@oRo�WR_C�ONFIG p.�%�c�_��IDL_CPU_kPC�PB�����` BH�eMIN��l�!�eGNR_I�O����`NP�T_SIM_DO��f{STAL_oSCRN�f �z�TPMODNTOqL<w{�QRTYxp�a	v@K0ENB<w��#�cOLNK 1q�� ������&�8��rMAS�TE�`�y`R�qSLAVE r��H D�uSRAMCACHEV�h�M1O_CFG���s���UO'@����CMT�_OP�P�b��Y�CL��ʅ�P_AS�G 1s�g�
 :�]�o��������� ɟ۟����#�5�G�\B�0�NUM���
��IP����RTRY_CN��ʅ8qG_UP����q��� ��׀��tT_ � 0aT��`RC�A_ACC 2u��+  L[T�� #Û0� 6�4� 69b8�qT:�0�" #�@J�<�PB j���BUF001 2�v�+= ��u^�u0�Ľ�н��ܽ�꽴��������+�7��E�Q�`�m��y崇崓崡�崭崹���Ӫ���������U����!��-��U9��H��T��b��Uo��|�ĉ�ĕ��U��İ�ļ��˅�Uׅ���򽳋������&�2޽��3����T��[�(YpT����Tǖ�  ���Tt�uT��]��L�  LW�����������������2����˿u0n(���� �������������� ��������$���,� ��4���<���D���L� ��T���\���d���l� ��t���|��҄��ы� ������������ �������������� ���������������� ����������А�� ��А����#�(�,� (�4�(�<�(�D���K����S�L =x[�e��c�e�k�W0 s���{� }у��ыѐ�А��/!xS���3���� ���Ҋ��Ҋ�Բ��ܲ ������������� ����"���$�2��� 4�B���D�R���T�b� ��d�r���t���� ���¢��²� ������������ ��������� ��"��!#�2�1 4�B�1D�R��!S�a \�r�d�r�at҂��� �Ғ���Ң�d���;2w�+ 4a\lU*�!� <� ��\�b�HIS��y�+� �:� 20�18-02-27�&�S/e/w/�'<�  ;�/�/�/�/�/^�-LY�3,(58/�%?7?I?[?m??�;���Q�/�?�?�#N�2,'1�?OO(O��H�ـ�X�!�0`=DMhMDiC�jL�=D�2fO�O�OLM����8�W�?�O�O�"<P�!�O�&TB:ZGp=D%xMD�=D|E�=Dhj��=D�=D��_ 2L���8�A�O�_ �_�_�&DB5PLB�TJ �@R�0HR�P_b_tYs�ڂ_ 2K��8�1�_�o�o�o8N�0S1!�?�o�'��o#5�&J�n�8��o�u��<B5P�emf�^o���%xR5P�n2ST�	'��/(/b�p�������<�5  Z��ҏ�����/ ?c�P�b�t������� �8��ٟ��?�?!�3�E��i�dD@d�L@qdT@d�\@t�d@d�lO+ -�L�@6ɟ�� �O�O���Z��%[ ���@Pd�HPt�,`d� |@d�<`d�hd�pPd� xPd��P8��_�_ݿ� ��]X�L@d�y�d�@P t�HPd�u�����\`�� qo�o������\�t��` t����t�I�[�I [�ߣߵ��iX���)� �p�����X��X� �	'��;�M��ߕ������ ������ )�;�)���q������������<������ �GYk�j�U� LB -U� \B� d@��yC� �@���=*< ]^'[�@R� HR�  ,byE� <b� Db� pR 	�� �R���// (/�]�����[c �/����/�/?��c .?@?	y^?p?�?p߂� �?�?�??I/��rO�,O>O��bO+�I_�CFG 2za�� H
Cycl�e Time��Busy��Idl�B�Dmiz_L�AUp�F��ARead�G�Dow_H�O���CCount>�A	Num �B�C��dKF]���,�S�DT_ISOLCw  a�� �P�gNJ23_DSP_ENB  }Z�e�POBPROC�S�E�S�SOG_�GROUP 1{�}[d�< ��GP?v%�odO?"�W_Jo�Q`o�o �o�oho�o�o�o���_�X�PIN_A�UTO�T�W�SPO�SRE�_�VKANJI_MASKiv�QzKARELMO�N |a�O_�y �o����)�gN�rv~B}a��R��A�K�fxuCL;_LApNUM�P���}pEYLOGG'ING}�f�����U�mPLANGUAG�E a����DEFAUL�T ��O�LGAy~Y��s �j$?�  8�@a�u��'�7  ���t�9��B�;���
c�(UT1:\9��� ������ ��͟ڟ����"�4��]�(���J�LN_DISP }[��L_o]o��OCTO�L֠�DzgP�QA���OGBOOK ����W��AW�W���N%V�H�Z�l�~����������CĹ��	
�Q�a�F���E��_BUFF {2�}[ ��S�?�i�o��G�� �������� ���	�6� -�?�l�c�u߇ߙ��������߮�7�DCS� ���R=����� �;(�Ed�v��|���IO 2�� �@��@gP� ��������+�=�O� c�s������������� ��';K]o����ER_ITMz^d!�� $ 6HZl~��� ����/ /2/D/�槱SEV}���.�TYPz^��/p�/�/S-bqRST����SCRN_FLg 2���0�D� D?V?h?z?�?�?�?�/�TP��z_�"�NGNAM�T�E��7UPS��GI� ���UA_LOA�D�PG %�:%�HA_1�?�]MA?XUALRM�����@��U
�B%A_PR*D� ��Q�@C�����Ot�wM��@�PP 2�� �"f	�/I_4_m_ X_�_�_�_�_�_�_�_ �_!ooEo0oio{o^o �o�o�o�o�o�o�o AS6wb�~ ������+�� O�:�s�V�h�����͏ �����'��K�.� @���l�����ɟ۟�� ���#���Y�D�}� h�������ׯ¯��ޯ �1��U�@�y���n�𯿚�ӿ|HDBGDEF ��58��O��_LDXDIS�A
@�;��MEMO�_AP@E ?�;
 ���]� oρϓϥϷ����τ@�ISC 1��9:�ƿ(�´�>����w�bߛ�
���_MS�TR �l-��S_CD 1�L͠�� ��1��U�@�y�d� v����������� �+�Q�<�u�`����� ����������; &_J�n��� ���%I4 Fj����� ��!//E/0/i/T/ �/x/�/�/�/�/�/? �//??S?>?c?�?t? �?�?�?�?�?�?O���MKCFG ���ݗ@XO�@LTAR�M_@B�WVB�*PB���O�D�@ME�TPU(�B�����NDPADCO�L�E��NCMNT6�O �EFN�@�O�G�� ���K^�C�VAc_mT�EPOSC�FW^PRPMl�O}YST�@1���� 4@@<#�
�QA�U�_g�_o oo[o=oOo�oso�o �o�o�o�o�o�o3�'iSq�ASING_CHK  _�$MODAQsC���TKVN�uDEV �	��	MC:>�|HSIZE(�@�ȣuTASK �%��%$1234?56789 D�V���wTRIG 1�.�� l��%�̡��C��ˏ����&�YP�����t�sEM_?INF 1�zG��`)AT&�FV0E0؏O�)�7�E0V1&A�3&B1&D2&�S0&C1S0=>>�)ATZO�����H��ϟ^�Ï����A��'��K�2�o��� 5���Y�k�}��� � ��$�[�H�Z��~�9� ������ؿ������� ӯ�V�a����ÿ�� k�u��ϡ�
���.�@� �d��)�;�MϾ�q� ��������<���`� r�Y��I�[���ߑ� ���&���J���n�)� 3��_����������� "�������|/�� ��������0�T�NITOR�4PG ?�{   �	EXEC1TC�2�3�4�Q5�g��7�8�9C�$�$ �$�$�$�$ �$�$�$�#U2	(2(2!(2-(U29(2E(2Q(2](U2i(2u(3	(3(�3��qR_GRP�_SV 1�$�� ([q�����&�޹�����+&���?g���}.�_D���]3ION_DB�B@��}A  ��@�x�?�2�x@V�A  N B��?�y-ud1��uO%O7OjAPL_NAME !;U�`@�!Def�ault Per�sonality� (from FsD)�1�ARR21� 1�L68L�@P`A�0
 d^R�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o�s2�ORodovo�o�o@�o�o�o�o�o�r<Ao 0BTfx�������?HBABD�
�B�ADP1� n���������ȏڏ� ���"�4�F�X�j�|� K�]���ğ֟���� �0�B�T�f�x����� ������������,� >�P�b�t����������ο���� �H�6 H�b GH\�AG70�0�C�U�ABd?�'�tφ�j� �϶�(��=J������8��!�$� �<� 2�D�V�t�zߘߺ�70Њ����AB�	`�&� �2�D��:��oA�Bd�v���? A�  ��BҏC�XI�0�@ � J`@�� @D�  ��?������?A@��AAA��6Ez  ��~?H;�	l�	� �@� 020��0E� ���� �? � �j�70�J��K ���J˷�J� ��J�4�JR�<�ܚ5�T���70@��S�@�;fA�6A��A?1UA��X������=�N��f������T;f���X�������*  ��  �5��>6 ����5Ȭ�N0�?����#�AA����5����`�������ҍ Vz0� (�0�� ��0���
��	�'� � (�I� �  y����:�ÈL?È=���d���� <E��� � �� ����=K����u�1��  '�0$�� @�!�p@�a�@j @ @!C5 KCF �F A B���CI�1�@�~������?�������_�_��@A@�%AAD ���/�/??>?)=�u�i!y5AC� :���  �x?��ff�Ϫ?�?N? !���?K��8A@O'J>�ל��� TFP^Hy9[�T�T���>����1�<�2�!<"7�<�L��<`N<D��<��,���O�?�����DB���?fff?� ?&�P��@T�Q?��`?Uȩ?X�(Q�p"Q� P
��\_��{_�G@��? �_�_�_�_�_�_oo�@oRo=ovo�EUF � eo�oao�oM_�oqY��o*�hHmN H�[��G� F��3l~i�� �������D� /��m�1���o�� ڏM����"�4��OI� [�����y�����֟����"q  ���� C@П5�̟Y�D�\ �c��j������ç�¬�q�BHF �R ���P��}�|� �@�Iܸ�@n��@��@: �@l��?٧]�� ��%��n�߱���=�=D��T��f���@�o�A�&{C/� �@�U|�
 +J�8��
H��>���=3H���_�� F�6��G��E�A5�F�ĮE���̿ް��fG���E��+E���EX���ް>�\�G�ZE��M�F�lD�
����i�Tύ�x� �Ϝ�����������/� �S�>�w�bߛ߆߫� �߼�������=�(� a�L�^������� ������9�$�]�H� ��l������������� ��#G2kV{ ������� 1.gR�v� ����	/�-// Q/</u/`/�/�/�/�/z��(��4��/�A��5�%3����/?�4 �{x ?2?��0+#L?�^?@2jbx?�?1?E�䴛|�@�; �9�?�?O�?,OL��%P�BP^Nm�z��O��/�O�O�O�O�I�0� �O�O'__7_]_H_�$`_r_�_�_�_�_�_@�Ol�&ooJo8lePo�Zo�o~o�o�o�o�a)�o�o8&\�jz  2 H��6�H��2�s\�b�B	���ݠB��
�A�@���֣@����5������y����������JTt���Q�9xv�
 ɏ� +�=�O�a�s����������͟ߟ����� ���H;���4��$MR_COM ��HH���z�3�x%% 2�34567890	1c�u� `������0��0ݡ�0�1�
���not sent *��1��WPET�ESTFECSA�LGRm`g�:�qd�(�灿�
8�kp�t@�4#�U�S�e�w���� 9UD1:�\mainten�ances.xm�l��ؿ  ����DEFAUL�TA�<�GRP 2=�G� �H����  �%1st� mechani�cal chec�k���1�t��|Å�lu;@H�����������ϒ2L�controller\�&�u�J�mt��v߈�0�߬߾��MS����2"8���0��lue�2�D�V�h�z���C߬�����3��)����"�4�F��C�U�geQ�. batteryJ����lu	����������
��Supply? greasoa1�3��H<�0RYlu�������z�^�cabl.E�1�
uJ\n ��Y��i���9/ /2/D/V/�Q �~/�<LH�/�B��/ �/�/	??j/??�/�/ �/s?�?�?�?�?�?0? OT?f?x?MO_OqO�O �O�?�O�OO�O>O_ %_7_I_[_�O_�_�O �__�_�_�_o!op_ Eo�_�_{o�_�o�o�o �o�o6oZoloA�o ew����o�  2�V+�=�O�a�s� �����͏��� �'�9���]�����Џ ⏷�ɟ۟���N�#� r�����W�}������� ů��8�J�\�1�C� U�g�y�ȯ�������� "���	��-�?ώ�c� u�Ŀ��追������� �T�)�xϊ�_߮σ� �ߧ߹������>�P� %�t�I�[�m����� ������:��!�3� E�W���{������ � ������l�A�� ����������� 2Vhz;as �����.@ /'/9/K/]/�n/�/ ��//�/�/�/?#? r/G?Y?�/}?�/�?�? �?�?�?8?O\?n?CO �?gOyO�O�O�O$K�2	 @�O�O�O&O_ ._@_R_d_v_�_�_�_ �_�_�_�_oo*o<o No`oro�o�o�o�o�ox�o�o  �\Aw?� �C _ =Oa�6)�����8*�**  6A8F}p��*��pN�`�r�����_O XC���Տ������ /�A������������ ��	�˟����c�u� ۟a�s���ϟY���ͯ ߯)�;�M��9�K�]������������6��$MR_HIST� 2�4E��� �
 \B$ 23�45678901P��ֿ�r�9�? k�}�4�f��?������ �ϲ��1�C����Z� �ߝ�T���x����߮� ���?�Q��u�,�� ��b���������)����M�_�����SK�CFMAP  �4E��~r�;�;�����ON?REL  ;��������EXCFE�NB��
�����F�NC��JOGO/VLIM��d��O ���KEY��R[_PAN��mi���RUNBnSFSPDTYP&<����SIGN�����T1MOTD�����_CE_GRP7 1�4E��� �@P;�=z�d �\�����/ 5/�Y//R/�/F/�/ �/�/�/�/???C? �/M?y?`?�?T?�?�?��?�?�;��QZ_E�DIT����TC�OM_CFG 1����	VOhOzO }
7A_ARC_��1	T_MN_oMODE��	UAP_CPL�O�NOCHECK� ?�� �� _&_8_J_\_n_ �_�_�_�_�_�_�_�_�o"o��NO_WA�IT_L�,GN�T?A����5;��ta_ERR!2�����|�o�o�op|���&Oe�@O�c���m| #��1�����W���v�n9�_��vB���<� v� ?�7��,��|�n�bPARAM�b]����t�?���8��1�C� =  G�`�r�z�T������� �����ҏ�,���7��^�p�����CU�M_RSPACE����}A͟ה�$ODRDSP�C��OFFSET_C�AR"@�O
�DIS���S_A�@AR�K�-IOPEN_FILE6��}A-F��PTION_I�Ocu��M_PR�G %��%$*�ǯٮj�WOV��'sv�
�;�t�  ��u$���$�	 �9�$���;���RG_D?SBL  ������j���RIEN�TTO��;�C�����A �UT__SIM_D�����r�V�LCT �~m)B�՝;�Z �_PEX�@9�(ķRAT�G d|(��UP ��
}�����Ϝς��Ͼ���$PALxb��~n��_POS_C�HW�5����p2 ��L68L@P>ݳ
 d��R� d�v߈ߚ߬߾����� ����*�<�N�`�r� �����9�2A��� ��� �2�D�V�h�z� ���s����������� "4FXj|�>��s��������bP �*<N`r �������/ /��J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?'/9/�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�}?V���O�M"Â�|q_  [_@_NW�M�M���_|_�_hW%��W�_�_ �_�_oo0oRo�P��0uo�l
t�T	`�_�ox�o�o�a:�o±��o0\�A��  Gy�'�Op�1�������� 6��b@ ��^���}p @D�C  �q�q�q|q?� ��q�D�  Ezx�s��;�	l�r�	 �@�� 0�@�A��p ��p� � � ����PH0#H���G�9G����G�	{Gkf��àWT��OP�b��PC�ᷰ��p&�D	�? D@ D�w?������  �O5��>���pú�������� B��Bp{�!�O��Oߔ��R ��&��q;��S�K��\��)��p�( W �p���Ј���_���	'� �� ĒI� ��  �Hp�[=����������� <�p� �� � �`�_�:��_��D�k��Nð�� C '԰��u��C��C���݀B�p�����ʯ� ���@�~2����.�?����G}±�nDp@� h��r�u ����}�����ڿŽ��#��ž� :���8�x?�faf__F�X�� �`��ϟ�ѱ8� ����>��8��qȺ��ƁP����q�s�tZ�>癙�<�@�<2��!<"7�<L���<`N<D��<��,(�e�t�Ɩs�N���Dp?f7ff?h�?&����@T싴�?��`?Uȩ?X��Ѽ	��ѩtȹ�u �ߖw���tw�L�7� p�[��������� ���$���H�3�l������e���a�HmN� H[��G� F���� >)bM�q�� ���o�	�[��� O��v����� o����*//N/9/r/]/P���"Ht�/� Cl/�/h/�/�-?���/???*?��Kç�s©-��H�E���O?<4�0�1�1@I���@�n�@��@�: @l��?�٧]�? ���%�n�������=�=D����?@��@��oA�&{C/� @�UO� �+J8���
H��>��=�3H��_@O �F�6�G���E�A5F�ğ�E��hOz@���fG��E���+E��E�X��Oz@>\�G��ZE�M�F?�lD�
�p�O �?_�O)__M_8_q_ \_�_�_�_�_�_�_�_ o�_7o"oGomoXo�o |o�o�o�o�o�o�o�o 3WB{f�� �������A� ,�e�P�b��������� �Ώ���=�(�a� L���p�����͟��ʟ ��'��K�6�o�Z� �����ɯ���د�@��5� �2�k�&B((A�4�o�(���<��X�3�ϩ����A4 �{��οA��0+#���ܲ�jb�&�1E����|��B�@ɀ�nϠ�ϒ��϶�)P`�P��-#�v�/�Y�D�}�h�A���ߊ��� ��������B$��� G�2�k�V��6���������e����,��0<�b�P�.)h�z������������
  �2 H�6FHY�;�'\�FB�!L�!y0BȎ0�0A@@�/n������/��'9�K]D��@�@�@E
 e����� /!/3/E/W/i/{/�/��/J� �������4�$PAR�AM_MENU �?@���  DE�FPULSEK�	WAITTMO{UT;RCV?� SHELL�_WRK.$CU�R_STYL0�B<OPTXX?P�TBm?g2C=?R_DECSN0�ž< �?�?�?O OO$OMO HOZOlO�O�O�O�O�O��!SSREL_IOD  <����E�USE_PROG %�*%�O>_�CCCR0�B��#QW�_HOST !F�*!VT�_KZT�]_�Sv_�Q�S�_J[_TIME2�FfU�� GDEBUG��@�+�CGINP_�FLMSKoCiT�RRoCgPGAp` 23l��kCHQoBh�TYPE�,�  �O�O1,>Py t������	� ��(�Q�L�^�p��� �������܏� �)� $�6�H�q�l�~������EeWORD ?	��+
 	RS�q`��PNS���Q4��JO�1��TyE�P��COL�����@��gTRACE�CTL 1�@�]�! ���������d�DT Q�@����D 7� ��ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�A�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������ï #5GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ Sew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q�G�ߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� ����������/ ASew���� ���+=O as������ �//'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�?��?�?�3�$PGT�RACELEN � �1  ����0��6_�UP ���e�A
@�1@��1_CFG �FE�3�1A�/D��3HOTHFM  ��TEBDEFS_PD �"L�1��0��0IN@T�RL �"MBA8�cE�APE_CON�FI@�E��A/DTI�0L�IDC�"M	XG�RP 1��G� l�1@�  �[��1A�?x�D P�DV�C2��WO��0dcD�Y�Y�A�@�&PTOEBFK��_ ´�S�_�[B �Pa�_�_�_$ooHo��1>'oY>a���fo�o�n�o =N?�=R�o�o �o�o%I4�oX��T���  Dz�s��0
��� -�S�>�w�b������� ���Ώ����=�(��a�o�)�1
V7�.10beta1�/D��B(��A�\)A�G��NQ��>�ײ�{����A����ff��A��p�AaG�?7�  ޑ@��OP�� o���+�=�/CAp��^b�D�u���𙯔�CQKNOW_M  _E*F
T�SV �9Y��E
���1� J�U�@�R���/B�]	S�M2S���0���	�AB�0����p���l�ٴ������@zA��.�`6�2�D̲�
QMR2S���TVi���_d�����MST2Q1 15�I��4�E�� ���^F��	��L�?� Q�cߕ߇ߙ��߽��� ����J�)�;��_�@q�������2��8ͱ�Ͻ0�< ���3P3
��.�@���4 ]�o�������5����������6'9���7Vhz���8������MAD��6 
F��OVL/D  K����PARNUM � �ˁ���SC-HN 
E
��8��3%UPD���UO/��_CMP_0���0@�0'*Eg$�ER_CHKu%`(Cٲ�&r/�+RS��ů
Q_MOP�/�%�_�/��_RES_G���K
���_d? W?�?{?�?�?�?�?�? O�?*OONOAO4&5	�1<A?sO&5\�O �O�O(3���O�O�O(3  _-_2_(3U M_l_ q_(3� �_�_�_(3� ��_�_�_(2V 1����1ͱ@`|���"THR_INR�0!��5d^fMA�SSko ZgMN�jo�cMON_QU?EUE ���ΦT0c� 4Nl U�!qN�f�h�cEND�a?yEXEu1 �BEp�o�cOPT�IO�g;�`PROGRAM %�j�%�`)o��bTA�SK_IPb~OCFG ��o��^�pDATA��� �@#�2صf�x� ������Y�ҏ������ŏ>�P�b�t�'�IWNFO���D���d 0�͟ߟ���'�9� K�]�o���������ɯ ۯ����#�5�������D� _I�q� DIT � �����>�tWERFL<xQc���RCALL_C?ONF Ƅ�����%�0�@��R���ݳKN�p?�� 0�ڶL�DBD 1��.�]���/���VLdp�%�7�I�[� m�ߑߣߵ������� ������&���J�\�n� �����A���� !����&�8�J�\� n��������������! ������2��Qc u�!������ ,>Pbt� �����// �7/I/[/��//� �/�/�/�/ ??$?6? H?Z?l?~?�?�}/�? ��?�/OO/OAO�? hO�?�/�O�O�O�O�O �O
__._@_R_d_v_ �?�_uO�_�_O�_o o'o�_No�Oro�o�o �o�o�o�o�o& 8J\7o��_�� )o���1o"��go X�j�|�������ď֏ �����0�c�f� ���9�����ϟ�O� ���M�>�P�b�t��� ������ί���� I�:��3�p������� ��ǿa��!��$�6� H�Z�l�~ϐϢϴ��� ������׿ �S�D�V� ɿw߉ߛ�ѿ��Y�� ��
��.�@�R�d�v� �������߽�� 9�*���K�]�o����� ��?�������& 8J\n���� ������C�1C Ug������ ��//0/B/T/f/ x/�/�/w�/��/�/ i?)?;?qb?�/� �?�?�?�?�?�?OO (O:OLO^OpO�/]?�O �/�Oy?�O�O_!_�O H_�O�?~_�_�_�_�_ �_�_�_o o2oDoVo �OzoU_so�o�O�o�o �o�o.a_Rdv �������� �*�<�`��o���� 	��ɏۏ���G 8�J�\�n��������� ȟڟ����C���F� y�j����������/� ��-��0�B�T�f� x���������ҿ��� )�����Pσ�qσ� �ϧ�A�������� (�:�L�^�p߂ߔߦ� �����߷� �3�$�6� ��W�i�{�Ϣ�9��� ������� �2�D�V� h�z��������ߝ��� �
��+=Oa�� ������ *<N`r�� ������#/#/ 5/G/�n/��/�/�/ �/�/�/�/?"?4?F? X?j?|?W/�?��?�? I/�?	OOQ/BO�?�/ xO�O�O�O�O�O�O�O __,_>_P_�?=O�_ �?�_YO�_�_�_oo_ (o�_mO^opo�o�o�o �o�o�o�o $6 i_Z5oS��_�� ����Ao2�D�V� h�z�������ԏ� ��
���@�sd�v� ���������y�'� �*�<�N�`�r����� ����̯ޯ�#�ݟ&� Y�J���k�}������ �џҿY�� ��,�>�P�b�tφ� �Ϫϼ������Ϳ� 9�:��[�m�ߑ��� ��O����� ��$�6� H�Z�l�~������ �������� �S�A�S� e�w������������ ��
.@Rdv �������� y�'9K��r	�� �����//&/ 8/J/\/n/�/�m�/ ��/��/??1?�/ X?�/��?�?�?�?�? �?�?OO0OBOTOfO �/�Oe?�O�O�/�O�O __�O>_q?b_t_�_ �_�_�_�_�_�_oo (o:oLo'_po�O�o�o _�o�o�o!_�oW_ HZl~���� ���� �SoV� �oz�)������я?� ����=.�@�R�d�v� ��������П���� 9�*��#�`������� ����Q�ޯ���&� 8�J�\�n��������� ȿڿ�ǯ�C�4�F� ��g�yϋ�����I��� ������0�B�T�f� xߊߜ߮������� )����;�M�_�q��� ��/����������� (�:�L�^�p������� �������� 3�!3 EW��~���� ��� 2DV hz�g����� Y//+/aR/�� �/�/�/�/�/�/�/? ?*?<?N?`?�M/�? ��?i/�?�?�?O? 8O�?}/nO�O�O�O�O �O�O�O�O_"_4_F_ y?j_EOc_�_�?�_�_ �_�_�_oQOBoTofo xo�o�o�o�o�o�o�o ,oP�_t� �_���o��7o (�:�L�^�p������� ��ʏ܏� �3�6� iZ�	�{�������� ؟o��� �2�D�V� h�z�������¯ԯ� �
���@�s�a�s� ����1�������� �*�<�N�`�rτϖ� �Ϻ��ϧ���#��&� ��G�Y�kߡ���)�׿ ���������"�4�F� X�j�|����ύ��� 	�����-�?�Q��� x���߮��������� ,>Pbt� ������� %7�^����� ���� //$/6/ H/Z/l/G�/��/�/ 9�/�/?A2?�/w h?z?�?�?�?�?�?�? �?
OO.O@Os/-?vO �/�OI?�O�O�O�O_O _�O]?N_`_r_�_�_ �_�_�_�_�_oo&o YOJo%_Co�o�O�o�o �o�oqo�o1_"4F Xj|����� ����o0�coT�f� �o�������oҏi� ��,�>�P�b�t��� ������Ο���͏��I�:��[�m������$PRCALL_�VER  ���T���W�ORK 2̰��� 
 \pG�����Q�( �� W�2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� ��������*�<�N� `�r߄ߖߨߺ����� ������� �R�0� �V�|�������� ������0�B�T�f� x��������������� ,>Pbt� ������ (:L^p��� `���� //$/6/ H/Z/l/~/�/�/�/�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O0�� �O_�0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�&_������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��t�ʿ���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������س��$PRGADJ� �ֵ��A�  *�? �4�7�d?��NS_�CFG �ֵ��?�  �Bz?�7�@7�<@5�?�k�%�k�������k�J�GRP� 2�X�'� 	_H  l����e�?z�A ?�ɻt$* / **:%7��*Fҷ`Է�� ��?�R�bt� ��$�� �:Lzp��� ����h//$/R/ H/Z/�/~/�/�/�/�/ @?�/�/*? ?2?�?V? h?�?�?�?O�?�?O �?
O�O.O@OnOdOvO �O�O�O�O�O�O\__ _F_<_N_�_r_�_�_ �_�_4o�_�_oo&o �oJo\o�o�o�o�o �o�o�o�ox"4b Xj������ֶ	 :�q�\��� ��	����叀�	���H�PREF ��X�7�7�
F�I�ORITY  �k�$�7���MPDSPON  ����v�UTb���K�I��ODUCT_ID� ����O=G��_TGLb�!����TOENT 1�����(!AF�_INE��2�=��!tcp=�e��!udT���!�icm|�����XuYQ��� �?�)� 2��7���,���X�?�|� c�u�����ֿ����� �0��T�f�*��Q��X�����ϻ�?�>W5H�,�2/<H���k������Az�,  �N���e�w߉߭��7���?�Q�/��PORT�_NUMb�7��m��_CART�REP��֬H�SK�STA�� �L�GS/�����z�7�Unothing��r���%��6�TEMP �����-�Z�_a_?seiban�� ��;�&�_�J���n� ������������% I4mX}�� �����3 0iT�x��� ��/�///S/>/ w/b/�/�/�/�/�/�/>��VERSI��&0 dis�abled ?SA�VE �Ě	�2670H755�(�/�?!�τ?�?���? 	�8��/�K	OR�e$OMO_OqO�O�J<L�?�O��F2]_� 1��o0P���u__�w0��URGE_ENB�����m�ǡWFKPDOb�7ү�W+�lT/����WRUP_DE?LAY ��_U�R_HOT %�T������_}UR_NORMAL�X̒�_<0o�WSEMIo5o|to.�QSKIP�C	ܹ��Cx�/�o�/�o �o�m�2 Vh z@������ ��
�@�R�d�*�t� ������Џ⏨��� �<�N�`�&���r��� ��̟��ܟ��&�8��J��U�$RBTI�F�	�RCVTMkOU���h��DCR�Cޗi ���aBcg
�BްB
W�A
<:���*F���m�cw�|����s�U?�3Pm�o�� <2�!<�"7�<L��<�`N<D��<���K��O�x��� R߮���ҿ������,�>�P�b�tϤ�RD�IO_TYPE � �Mj���EFP�OS1 1�N9��x�?��Rg� �� D��?h�ߌ�'߉��� ]��߁�
��.�@��� ��'��s��G���k� �����*���N���r� �����C�U������� ��8��\��Y� -�Q�u�����XC|��OS/2 1�[��3�m�i/���3 1���/�/n/|�/%/S4 1�</�N/`/�/??<?�/S5 1��/�/�//?�?�?�?O?S6 1�f?x?�?�?BO-OfO>�?S7 1��?O�OYO�O�O�OyOS8 1�O�O�O�Ol_�W_�__SMASK 1�� ���_�VN�WXNO���Vo<c��MOTEo����T3a_CFG ��:m�Qa��PL_�RANG6ar�taO�WER 鮥��`�fSM_DRY�PRG %�Z%�7_�o�eTART ��n�jUME_�PRO�o�oIT_�EXEC_ENB�  _�z�GSP�D"pdplx��{vTD�B��zRM��xI_AIRPUR}`� �_��]MT_��PT�`8k~�h�O�BOT_ISOL�C�^iffeD�N�AME �z�8��OB_ORD_NUM ?�h��qH755  ��֏����h�PC_TIME�v�xh�S232�Sb1뮩`�L�TEACH PE�NDAN��OWh�W�6_!Mai�ntenance_ Cons��f��"��No UseW���y�ן��������2�NPO��`�a(��/�CH_L%p��3�R	��l�!OUD1:ǯn�R�P�VAIL�������&�.aSPACE1w 2���k�@nbO�E�USP�nb��|���< �@�?�﫫�﯋��� ٿ��?�Q�c�u�'� �������ϑ������ *u.q'�C�U�g�y��� �Ͽϵ��ߕ������ !�;�Q�c�u߇�9�� ����������;� M�_�q��5������ ��������+I�[� m������������ �$�EWi{ �?�����  //5/Sew�;/ ���/��/�/?�/ ?O/a/s/�/�/I?�/ �/�?�?�??*OO?O ]?o?�?�?EO�?�?�O 2O�O_&_�O;_t�&�2+�� =�sO�O �OI_�O�O�_6_�_&oGoo\o]_3p_�_�_ �_�_jo�_oWo�o Gh?}~o4�o�o �o�o�o��o/2�x@�h���`����5� �������P�S����3�����������6 ӏ���	��͟?�q� t���T���˯����7����*�<��`� ����ۯu�˿�ÿ��8�'�9�K�]�� ��������������ϼ"�#�G �9�� �ZD
�� r�  9ţߵ��� �������;�v�.�]� ;�Z�ߍ�]Ad���� �����������"�4� *�<�N�?�|������� ��6���&8J @�R�d�v������� ��V"4FXj�`r���� `� @`@%k� /��	O!y�`/ r/xR*S/�/�/�/�/ �/�/!?3?�/??K? �?O?a?s?�?�?�?O �?�?AOSOO'O9OkO��OoO}
1/_a[_MODE  9ɼy�VS �9��O����-/V_�_��Z	�_�_�dCWO�RK_AD(\�
��4��aR  �9�F�?`�_)`_I�NTVAL(P�Đ�A�QfOPTION�`f ke�pV_�DATA_GRPg 2�D�D� P�_�o�_�o�i�O 	?-cQ�u� ������)�� M�;�]���q�����ˏ ���ݏ����I�7� m�[��������ş� ٟ���3�!�W�E�g� i�{�����կï��� ��-�S�A�w�e��� ������Ͽѿ��� =�+�a�Oυ�sϕϻ������/Q�$SAF�_DO_PULS�`0P�a�	���CAN_TIM'Q��e��R ����`��P^5P�����S�a�Rg�}QY�� �o�ߣߵ������� z��!�3�E�W�i�sX+��2��Y���d����bW�t� Cn����	�r����� �`��_; "  T>`/��l�~�����T D������������  2DVhz�������c_yU���0B�	!|iў;�ot�zTpbe 
�t��Di�Tiђ[  � ��}Q7Q i�a�Q����
// ./@/R/d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�Oq�,��O �O�O__'_9_K_]_ �O��_�_�_�_�_�_��_oo+o0am_r0 *�)��|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L��Op��� ������ʟܟ� �� }_6�H�Z�l�~����� ��Ư1o_eio��� *�<�N�`�r������� ��̿ڹ����#�5� G�Y�k�}Ϗϡϳ��� ��������1�C�U� g�yߋߝ߯����ߨ�������-�?�Q� c�u���������@����)�;�I��R������rb�x�N	1234�5678�h!?B!ܺ��s�|��% 7I[m�� ����&8 J\n����� ���/ /2/D/V/ h/z/�/�/�/�/�/�/ �/
??��R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO1?�O �O�O�O�O�O__&_ 8_J_\_n_�_�_�_�_ �_�O�_�_o"o4oFo Xojo|o�o�o�o�o�o �o�o�_BTf x������� ��,�>�P�b�t�3 ������Ώ����� (�:�L�^�p������� ��ʟ��� ��$�6� H�Z�l�~�������Ư@د���� �q���B�T��y�������Cz  Bp��_   ���2r�_ } ��
����  	�q�2@:�!�3�E�W�g���h��ϭϿ������� ��+�=�O�a�s߅� �ߩ߻��������� '�9�K�]�o���� �����������#�5�@G�Y�k�}�����h�t�ܲ<�� ��~�  ������Ƕ����t � Ѱ	 ǵ�$�SCR_GRP �1��@��# � ��� ׵	 _g�o �yi���ٵ�	���p�������6�C���}͆�$���LR �Mate 200�iD 56789�0�LRM] 	LR2D d~s�
1234c��v�g��첶 oǶ^�^�ù��}
��	�/'/�9/K/]/Ǵ��#H�o �s^�/���/�/�/�!�s���/"?�/F?��7?��hZ��,�	B���Ƒ?ȏ2�4�AѰ�?  1@��5�@��0�?# ?�5�2H��O��:�F@ F�`2B:O1?^OIO�OmO �O�O�O�O�O _�=�1��2+__(_:_LTB� Z_�O�_�_�_�_�_�_ �_o	oBo-ofoQo�o�|Ϛj��g�o׷����os��1@>'�1U�@�0O���ew���9��ǴA�0�f�u�/��%�p���s�  ��$�2� �G�S�$e�4�f���
����������o�̏�7ECLVL  s������rA���*SYSTEM*��V9.1035� P�7/19/2�017 A ����>�e�SERV�ENT_T  � $ $S_NAME !���PORT����R�OTO�� s�_S[PD{�(� ����TRQ  { 
��AXIS��9���� 2�`���DETAIL_ � l $D�ATETI����E�RR_COD�I�MP_VELϰ� 	�TOQ �A�NGLES �DI�Sz�,���G��%$�LIN�����R;EC�� ,��ʕ��$�MRAn� �2 d��ID�X��i��� �f�$OVER_OLIMI��Đ	g��OCCUR�� � �COUN�TER�� �SFZN_CFG��� 4 $EN7ABL�ST ����FLAG��DEBuU$�R9� g����D �� � 
�$MIN_OVRD��$Iy�5�Y�<Q�b�FACE��Z��SAFy�MIXE�D��b�B�Y�ROBކ�$NE��PP���h�HELL��	 5$J���BAS�RSR_��  $NUsM_�� � �1U���2�3�4��5�6�7�8�U��ROO��\�C�Oy�ONLY�`$USE_AB����ACKENB����IN��T_C�HK��OP_SEsL_���_PU����M_�OU��PNS����ԳV�����M�TPFWD_�KAR����RE���$OPTIO=N6�$QUE�ɝ��D�YͲ$CST?OPI_AL��Գ�EX����j��XT���M1��2��MAn^�STY��SO���NB��DI��TRqI$�b��INIz�9M����NRQ�և��END��$KEYSWITCH�����k�HE�BE�ATMM�PERM'_LE�%�E�L�U�F���S��D_O_HOMy�Oͱ��EFP����%�А�ST*��Ce�OM|�n�OV_MS�����ET_IOCM�N��rװ�;�ճH}K{�
 D �f��SU�`�MP����PO��$FO{RC�WARN��OM�� �0�$FUNC���UL����AR��h�2g�E3g�4\�;���O*��LM�w���UNLiO�����ED����SNPX_�AS� 0�A�DD4�6�$SI}Z�$VARU��MULTIP�����l�AM� �� $�����	�����C�IF'RIF����SJ�\���9 NF��ODBUS_AD���	��;���|� �� ��6�TE��$DUMMY8��SGL�TA��  &����`<� � STMTj��PSEG��BW<e��SHOW���BANTPOF4b�9�10X�ѭh�VCy�GF� � $PC����x�£$FBI�P�SEPr�A���tDz~E�� ���A00?��p���z��������5��6�7�8�9
�A�B�[���� �F�b�(�U1�1�1
)1)�1$)^��(>)1K)1�X)1e)1r)1)1��)1�)2�2�2��2�2
)2)2�$)21)2>)2K)2�X)2e)2r)2)2��)2�)3�3�3��3�3
)3)3�$)31)3>)3K)3�X)3e)3r)3)3��)3�)4�4�4��4�4
)4)4�$)41)4>)4K)4�X)4e)4r)4)4��)4�)5�5�5��5�5
)5)5�$)51)5>)5K)5�X)5e)5r)5)5��)5�)6�6�6��6�6
)6)6�$)61)6>)6K)6�X)6e)6r)6)6��)6�)7�7�7��7�7
)7)7�$)71)7>)7K)7�X)7e)7r)7)7��)7�$f�VPI�U�� ��V���
t�{���$7TORS�CMX�"��M��R��ǰ �Q_ҠRx�.�ϑ%� �h��YSLS�|� � ����x��(���x�؄�VALU����֨��FɁIgD_L��9�HI4��I;�$FILE_���d���$��ĆS�A�� h ���VE_BLCK�Mӝ����D_CPU�������g�y���ŁV���R ? � PWԠ��lp �LAS����-�&�RUN_FLG?��C�&��F�d��d�&�H��2���|&����TBC2C� �� ��F����චk�Ծ���TDCF�#�עQ�b�ҧCTH�� ����R��~��ESERVE��-���-�3������� X -$X�LEN��e���X�Ɛ�RAIд�ȀW_����1X�Q�2��MIO����S� ��I�����]�ǹ��X�ܻDE<�LACE�ⱃ�CC��]�_MA����%���%�TCV,�M���T��N�m�c�@�곖�����J���M���J���)����d�2�Ћహ���*�JK�V�K������N�
�J�c-��JJ!�JJ)�AAL�O�!�O��I�4J�5
���N1�t̀�?�)���LŰ_�����CF�� =`��GROU����қN��C1��R�EQUIR��E�BUHT���$T�2�U��֞��� \��APP�R�CL��
$O�PENN�CLOSD��_�S��s��
��. �5�M�*�8�(���_MG`����C�����'���B{RK��NOLD��>2RTMO_���$���J��PQ�� !��)��m��v��%6>�7>������� ��l����!Ѭ�PATH ������񄸽� �9��xSCAB��lO��INW�UC˰�� C�UM Y������'=�3�B
�!�B
N�B PAYL�OA��J2LY�R'_ANߡ�L��	��}	���R_F2�LSHR'��LO���4�4ACRL_��ur(�H���$H���5FLEXQ��:��J�� P;⳯�ů,�>���RW� :d�v������y�)���������F1 �,%@'��ǿٿ����p"E�+�=�O�a� sυϗϩ�G8d4���� �T v8���������	T�7E1X��N1ճ$ �(�E�(�*�<�N� R�[�I�m�v߈ߚ߬�sSTQ�� ���`�������Z�ATY&��EL� k�+S
�J��JE��C3TRT!TNt�'V���HAND_VB⯂Q���  $��0F2�����S�W����!� $$M� �阀���X@���\
0�U,�fA@� z ��?�#i��A���
��A��A��.`��ϐ���D��D��P��G9��iST���a���aN��DYE�L���d 6e� Y�����| כ4 �0�PF�O��X�a�j�s�|���R�J��"�P+R���r�v<���qASYM����	���!0�_��� /���X 9K]o�J�9���
�����	f$_VI�S�����V_UCNI'��>C�J� 5�cu5��9��F�j� ���9�,���3IBJ�P��H��@�#�R�d�D	I����O
�����C�$ N@=bI �A =�47�Z E�E�] l����� � % �[ �QME�!�@h`���G�T��PT�� �@�������Dc�ȍ�����T���� �$DUMMY1�N�$PS_W RYF ��$���7FLA��YP�3�����$GLB_T �P ����l�� XQ�d�& X;��ג�SuT�!�SBR���M21_VK2T$_SV_ER� Or�L^�v�CL2�^�A� �O:��GL��EWοq' 4�В�$Y�bZ�bW�����r�SAa�  ��]U��( �0N۰ޣ�$GIhP}=$�� '摤�ڰ�q) L����q��}$Fq�E�NE+AR� N^#FKɦ �TANC^" ��JOG /� �*�P$JOIN�T�1	@���MSE]T�q+  ��E1��!�@S�B�@��@�q_,� `PU�!�?��LOCK_�FO� �Q�BGL�V[SGL��TES�T_XMQ��EM�P��K2�0���c$U����02(��ڳ?�)
ҳP��?�'�`�CE���`� $�KAR1M�TP�DRA��}�t�VE�C���x�IU?�*�D�HE��TOOL� #��V$RE��I�S3���6a�T ASCH���+��O��L��Ҥ29ۢ��IA��  @$RAI�L_BOXE�1ރ�ROBO�?�~��HOWWAR=x/����ROLM� U�A��f��A�H ���O_F�@! �	���ѿq-�΋�R
��O�.�� ����Y�R��OU��/F��;�'G�1RQ��$PIP�N�0������f ?Ѡ�CORDED�������@�OG� 0 D �OBca5S��R��A�̣�A�q�7QSYSA�ADR6Q琈��TCH�P 1 M,�0EN�mA���_�����AE�C_��VWVAc�2� � �Ч� �P�REV_RTpq�$EDIT��VSHWR�AJ� �"J����Dr��)~>A$HEAD��h��C ����KE���ƠCPSPDZJKMP^�L��PR� F"�3I�b��I�5S6RC|PNE��7Q�rWTICK #*�M�k��HN@�4� @K��Eb_GqP��nSTY����LO2�㰱����p5 t 
��G���%$����=J�S,@!$+��0w���4��P��SQU�w�%���TERC܌��r�TS�D6 �V��G�0�GC1Ī�G�O����b IZh����ߡPR3�0�"���PU�A%g_DOP­�XS���K��AXI> y�D�URP�#7R6�� �l��QP_��~�ET�"P��Z��u=Fd�w>A�a�Ӥ���NA!�R�T7l��YB �Z�%�V9b�%g�# i�#/i@5Qg@5ag@5 qfR5l=�iR5�<�rp9B�;~=C�=j�|���ܠ��qSSC� 78 h��DS� ~�fҠSP1�lEAT_`�b !� �ϢAD�DRES��B��S�HIF�C6�_2C�H6Ph�I9��A��TU9�I�Q 9>��CUSTO�$q�+TV��I%�:����A#�p
�
�q�A,$B�; \H�����=\��KRC��c��"Z��|�KQ�TXSCREEC��<��YTINA��
��T�����!�B�p= T�y�"~� x�U��VL!}�L"�T��RRO:pe�}�T �Q�V���UE�> ���p���S��~�RSyM� B'UNEX���Ua�S_Գuf$� eaxi�g$��!C��Qb��T 2=�UE¼t?+����f GM�T}�LW�[!e�O~���BBL_��9W��B�@ �=r5Oα!rLE�B,sx5��B+tRIGH5s�BRD���ACKG9R��]uTEXn ^u>YqWIDTH� �U������ �U�I��EY�@qA Ad��z T�!�!BACK��u���k�FO*��wLA-B*1?(k�I����$UR;�����p�q�Ha B 8�̑e�_B�B3�r�R�������ڢ�� �O��ApC� ��VpU�Ap��R��`�LUM8��c&�@ERV����PO��tDi�� G�E�6�� ��)K LIPӅ�"E�1A)��@AA��QA������5��6��7��8������
 O�_TѦ����Sv�C�qUSR��OE <H�q�U ���C �FO�@ �PR�I�!m�o�ҐTR�IP�m�UN�#�F��b�D%�G�C%�p7�} w qG.���!G JaTy�A�A)�OS���>�R� b���qH���³ɾe��7�UہqIn����cۂ N�OFF�pJF����O�� 1Hh��ޤ�I��GUx�P���!�A+��qS�UB���`SRT�g��$K�d����O9R��q�RAU� r��T�������S��A �L HK�SHA�DOW` �ӿ�_UNSCA�ӿ��t̳�DGD�ѵ��V�C"0G��aM� �B�nF�΂����C�� �DRI5V&�!_V� C��� T�D~�MY_UBY}�(�De�na���P0���ѽ�P�_հ��L%+BMv(q$� DEY���EXp)c��t _M�Ux X(q�j`US |��͐�еPt��@�bu�G�0PACIN�kRG1 K�b��̣bҋ�bҝc�REH��A��r�bҝ��N ��TARGBh�P"R�����RU����O�pz�M!�qQ�	l�<!RE�SWZГ_A[�p� OD���AA�@��"En��U0J�q�p�HK5P� 3��!���Pd�EA� n�W�OR5���MRC]V�aQ �̀OAM5�C#S	��ޣ����REFw���� 
ཀ�#�Т����������%���Z�_RCo�[���z0Sk��t���}�0��dR �@�p�u���y���OU��� (� SM�� A2�0$�PaP � OC A��K_ SUL#PPf��COI`J�Q� NT���PE��O b�O��O L��x`��xb������>�S� ,C�!zB@ CCACHLO������	c!��@�C_LIMI�CFRTX0���$HO5���� C'OMM>�QbO?pG`��� ρ��H@VP��$���_��ZFЏl�WA MP�WFAIG`�� �AD���IMRE��"�GPW`��� ��ASYNBUF�VRTD6%B$�6psOL�@D_ƣ^%uW��P�0ETU���� Q8�&%ECCU��VEM~���"VIRC�V%>#Pb>B!_DELA��W�X�鐪�AGR)R�GXYZ�`c�W���3�q� T���IM��!U%��dT�B�qL#AS�pq�_� !���U���S �N��4��LEXE�V��S����A�FL2ZpI��(#FI` �7Ű�8��a���!�0
��W���:�􂔊�\��,pORDƑȧѨ�C��pX�P��T��b��O�p���sSFxp9cY  �P��O�UR����S�M�Z����$A3DJR@����U�[��oG2�LIN��Q`�XVR�\|Z2�`T_OVR�2���ZABC^�]��3R"CwQ�  ��Z(��^����$L�t��r��ZMPCEF^�_�B�P��Rn��LNKr
�Q	�_�` �̀Tn�^�TCMCMT�C��CART_�Q-�P<����$J�S�TD�Rbg	�e	��/�UX!1�UUXE�@f!1e8deca�Ia[iIakf�ZZU�a �KuT��aY�PD�� b.�R�ő0HEOtРpGr�W�q��a>��c � |D��QPWpEAK׈�K�_SHIF��HR�VF����<r(PC Xp�R�Q!}@8�Wq�P�V�IstD�xTRWACE�Vt��a�SPHERq�d� ,
 �h�o�i��f��aFA/����?����t�HOTSTA����MIPOWER�FL ����8�WFDO� �� �q����1 ������/� L{!��_EIPH������j!AF�n ��Əυ!FTd�������!���@��	�f�!R�{ MAINg�I��@U���y�n0��H������!TPn �����d�J�!
PML�o@XYK���e9�����d���f���!/RDM�0V㯰��gѯ.�!R90d/���h�z�!
{��T����ii�ƿ!�RL3 Cǿ�8|���!ROS���9��4�^�!
C�E�MTQ_ϳ�k,MϪ�!	s�Cq�ϲ��l����!s�W#AS���ϴ�m��B�;!s�USBC߱�n1ߎ�-����ߑ� �� ���$���H��l���x�I�pKL ?�%�� (%S�VC 1s���2����� 3���� 4��� 53�8� 6�[�`� 7���� 8H���� 9������ E� ���(����P ����x��%����M� ���u������� ��@����h��� ��>���f��� /��0/���X/�� �/��.�/��V�/ ��~�/��x��� ���C?�?��?�?�? �?�?�?�?OO@ORO =OvOaO�O�O�O�O�O �O�O__<_'_`_K_ �_o_�_�_�_�_�_o �_&ooJo5o\o�oko �o�o�o�o�o�o" F1jU�y�������~�_D�EV ����UT1:�4���&�GRP 2���O0��bx 	� 
 ,v����O2{�����܏ ÏՏ���6��Z�l� S���w���Ɵ���џ � �w�D���h�z�a� ����¯ԯ����߯� ��R�9�v�]����� ��п'�ſϽ�*�� N�`�Gτ�kϨϺϡ� ��������8��\� C�Uߒ�鿶��߯��� �����	�F�-�j�Q� ������������� ��B�T���x�/��� ������������, P7I�m�� ���[��:� ^E��{��� ��/�6/H///l/ S/�/w/�/�/�/�/ �/ ??D?+?=?z?a? �?�?�?�?�?�?�?O .OORO9OvO�O�/�O cO�O�O�O_�O*_<_ #_`_G_�_k_}_�_�_ �_�_oo�_8o�O-o no%o�oyo�o�o�o�o �o"	F-j| c������J�d ��	�1���U�@�y�d�����%�x��яQc���� �������(��L� :�p�~������f�П ��������N��� u���>�����̯��� ޯ �V�|�M���&��� n�����ȿ���.�� R�ܿF�ؿV�|�jϠ� �������*ϴ��� B�0�R�x�fߜ����� ߌ�������>�,� N�t�ߛ���d���� ������:�|�a�s� *�L�&����������� T�9x�lZ| ~����,P �D2hVxz� ��(�/
/@/ ./d/R/t/���/ / �/�/�/??<?*?`? �/�?�/P?�?L?�?�? �?OO8Oz?_O�?(O �O�O�O�O�O�O�O_ RO7_vO _j_X_�_|_ �_�_�_�_*_oN_�_ Bo0ofoTo�oxo�o�_ �o�o�o�o�o>, bP��o��ov� ����:�(�^�� ���N�����܏ʏ� � �6�x�]���&��� ~�����؟Ɵ�>�d� 5�t��h�V���z��� ��ԯ���:�į.��� >�d�R���v����ӿ ������*��:�`� Nτ�ƿ���t����� ���&��6�\ߞσ� ��L߶ߤ��������� "�d�I�[��4��|� ���������<�!�`� ��T�B�d�f�x����� �����8���,P >`bt���� ��(L:\ ������� / �$//H/�o/�8/ �/4/�/�/�/�/�/ ? b/G?�/?z?h?�?�? �?�?�?�?:?O^?�? RO@OvOdO�O�O�O�O O�O6O�O*__N_<_ r_`_�_�O�_�_�_�_ �_�_&ooJo8ono�_ �o�_^o�o�o�o�o�o "F�om�o6� �������` E���x�f������� ��Џ&�L��\���P� >�t�b���������� "������&�L�:�p� ^���֟�������ܯ � �"�H�6�l����� ү\�ƿ���ؿ��� �Dφ�kϪ�4Ϟό� �ϰ�����
�L�1�C� �����dߚ߈߾߬� ��$�	�H���<�*�L� N�`�������� � ����8�&�H�J�\� ������������ ��4"D������� j�����0 rW� ��� ���/J//n� b/P/�/t/�/�/�/�/ "/?F/�/:?(?^?L? �?p?�?�?�/�??�? O O6O$OZOHO~O�? �O�OnO�OjO�O_�O 2_ _V_�O}_�OF_�_ �_�_�_�_
o�_.op_ Uo�_o�ovo�o�o�o �o�oHo-lo�o` N�r���4 �D�8�&�\�J��� n����ˏ
������� �4�"�X�F�|����� �l�֟ğ���
�0� �T���{���D����� ү������,�n�S� �����t�����ο�� �4��+���޿L� ��pϦϔ������0� ��$��4�6�H�~�l� ������ߒ����� � �0�2�D�z�ߡ��� j����������
�,� ���y���R������� ������Z�?~� r������ 2V�J8n\ ~���
�.� "//F/4/j/X/z/�/ ��//�/�/�/?? B?0?f?�/�?�?V?x? R?�?�?�?OO>O�? eO�?.O�O�O�O�O�O �O�O_XO=_|O_p_ ^_�_�_�_�_�_�_0_ oT_�_Ho6oloZo�o ~o�o�_o�o,o�o  D2hV��o� �o|�x��
�@� .�d�����T����� �Џ���<�~�c� ��,���������ޟ̟ ��V�;�z��n�\� ��������گ��� ʯ�Ư4�j�X���|� ����ٿ������� �0�f�Tϊ�̿��� z����������,� bߤω���R߼ߪ��� ������jߐ�a�� :��������� � B�'�f���Z���j��� ~����������>��� 2 VDf�z� ����
�. R@b����x ��/�*//N/� u/�/>/`/:/�/�/�/ ?�/&?h/M?�/?�? n?�?�?�?�?�?�?@? %Od?�?XOFO|OjO�O �O�O�OO�O<O�O0_ _T_B_x_f_�_�O_ �__�_o�_,ooPo >oto�_�o�_do�o`o �o�o(L�os �o<����� � �$�fK���~�l� ����Ə��֏��>�#� b��V�D�z�h����� ������ԟ��� R�@�v�d���ܟ�� ����$SERV_MAIL  
�� ���OUTP�UT����@�RV 2v��  � (��xЯ\��SAVE���TOP10 2}6� d � ��ο����(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z�`�����YPy���FZN_CFGw ����%�j���GRP �2�燱 ,B�   A:�D;� B;��  �B4��RB2�1i�HELL��!	����I�J����>��%RSR���� ������"F1j Ug�������0�  �>�%0^p>|���x��)�uF2�d�v�e�HK 1
s� �$//1/C/l/ g/y/�/�/�/�/�/�/ �/	??D???Q?c?_�?OMM s��?�d�FTOV_EN�B��>���HOW_?REG_UI�?��IMIOFWDL�0�>=�BWAIT�2��0F��6�=�-ITIM�5��gOVA��>OA_UNIT�3�F���LC�0TRY�7����MON_ALIAS ?e�9E�he��"_4_F_ X_fZ_�_�_�_�_j_ �_�_oo+o�_Ooao so�o�oBo�o�o�o�o �o'9K]n ����t��� #�5��Y�k�}����� L�ŏ׏������1� C�U�g���������� ӟ~���	��-�?�� c�u�������V�ϯ� �����;�M�_�q� �������˿ݿ��� �%�7�I���m�ϑ� �ϵ�`�������ߺ� 3�E�W�i�{�&ߟ߱� �����ߒ���/�A� S���w����X�� ��������=�O�a� s���0����������� ��'9K]� ���b��� #�GYk}�: ������/1/ C/U/ /f/�/�/�/�/ l/�/�/	??-?�/Q? c?u?�?�?D?�?�?�? �?O�?)O;OMO_O
O �O�O�O�O�OvO�O_�_%_7_�C�$SM�ON_DEFPR�OG &����aQ &�*SYSTEM�*>_�W 	MWR�ECALL ?}�aY ( �}1�copy md:�prog_1.t�p virt:\�temp\=>1�92.168.1�.103:808;0 �Q868�_o�o)l}8�Rfrs�:orderfi�l.dat�Umpback�_�Quo�o��o,m/�Tb:*.*Rodomo�o"5d3x=d:\�oGp�o��Q�o��� }4=uaEW�Y����,mtpdisc 0��P��}������4etpconn 0 ^�X�j��� ��2oDo�ohoy��� ���o�o]��o��	�� .@�du��������O��t�����
�xyzrate 61ف˯ݯ﯀���䤿7�=�]�960 ؀]�o� ��$�7�˾ ڿ�}Ϗϡϴ�F�X� j�����2�D�͟λ u߇ߙ߬���Y�Ѹm� ���"�5���Z�ֳ�� ���﹯J�\�ٰr� ��'�:��������ȓ���8����U12884 ]�o� $7�11ō����z��1�2�_�_Np %��� J� ���7�HZl��/!/��Ƹ��07:798�P���/�/ �/7Ҽ_�M-p/?? %?8�J���Q)v?�?�? �߿�Z?R'm?�?O"O�545=?O8�/7:3�22�P�?�O�O*O-=F*.dQOcMkO�O _ _�E��O�O�O}_ �_�_4/F.nR\_n_�_ o#o�/�/�_�P�_�o �o�o7?I?�?jF�o �?�?�o�Y�o� �6�I�[�hHq�� &�����ldu����� �o�o�o^�t������<׏`򏃟���� ��$SNPX_A�SG 2����ȑ� �P��'%R�[1]@�����?���%���C�&� 8�y�\�������ӯ�� ȯ	���?�"�c�F� X���|���Ͽ���ֿ �)��3�_�Bσ�f� xϹϜ���������� �I�,�S��bߣ߆� ���߼������3�� (�i�L�s������ �������/��S�6� H���l����������� ����#O2sV h������ �9CoR�v ������#// /Y/</c/�/r/�/�/ �/�/�/�/??C?&? 8?y?\?�?�?�?�?�? �?	O�?O?O"OcOFO XO�O|O�O�O�O�O�O �O)__3___B_�_f_ x_�_�_�_�_�_o�_ oIo,oSoobo�o�o �o�o�o�o�o3 (iLs���� ����/��S�6��H���l���������PARAM ȕ�ґ �	��ÊP3�7�È�����OFT_K�B_CFG  � �Ε��OPIN_�SIM  ț��l�~������RV�NORDY_DO�  �A���QSTP_DSBU������ـSR �X� � &>�TYLE1��;�� �Y�ـTOP_?ON_ERR��ׂ~[�PTN X�����Cx�RING_PRMe��ȒVCNT_GP� 2W���x 	���֯���3���VD��RP 1	��$���n� ��������ݿڿ��� �"�4�F�X�j�|ϣ� �ϲ����������� 0�B�i�f�xߊߜ߮� ���������/�,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZ�~ �������  GDVhz�� ����/
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8O_O\OnO �O�O�O�O�O�O�O�O %_"_4_F_X_j_|_�_ �_�_�_�_�_�_oo�0oBoL�PRG_CoOUNT6�玢NgiENB��ieM�c�8��o_UPD 1}�T  
Wo  ��o�o72DV z������ �
��.�W�R�d�v� ������������ /�*�<�N�w�r����� ����̟ޟ���&� O�J�\�n��������� ߯گ���'�"�4�F� o�j�|�������Ŀֿ ������G�B�T�f� �ϊϜϮ��������� ��,�>�g�b�t߆� �ߪ߼��������� ?�:�L�^����`l�_INFO 1,�i�` �U`��������
�?���@Cz=��%���{���A�漸n ����³�vB���k`YSDEBUG�x`�`��d�i��S�P_PASSxe�B?��LOG ��e�a  r��M���  ��a���UD1:\x������_MPC����eI[�ay ��a)SAV ����a������SV}�TEM_TIME 1��]�` 0�`�����{�SK?MEM  �e�a�� %`r�X|�`�	�N� @��"��q��`�`��� ��/ �`)�� �@�?/Q/c/�   f-���23 ��/u( &"�/�/�/�,��/?0?B?�T?f?x?�?�?�?Hle �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O��O__&_8_�aT1?SVGUNS�`ye�'�e�MPASK_OPTIONx`��e�a�amQ_DI���o�UBC2_GRP 2;�c��_�6"0C��SA\BC?CFG �[�c �"k8m� Qo	�uo`o�o�o�o�o �o�o�o;&_ J\������ ��%�7�"�[�F�� j��������ʏ���� ����E�0�i�T��� ���T����۟ɟ�� �#��G�5�W�Y�k� ����ů���ׯ��� �C�1�g�U���y��� ������ӿ	��ڀ� /�M�_�q�ￕσϥ� �Ϲ�������7�%� [�I��mߏߑߣ��� ������!��E�3�U� {�i���������� �����A�/�e��}� ��������O����� +OasA�� ������9 ']K�o��� ����#//G/5/ W/Y/k/�/�/�/{��/ �/??1?�/U?C?e? �?y?�?�?�?�?�?�? O	O?O-OOOQOcO�O �O�O�O�O�O_�O_ ;_)___M_�_q_�_�_ �_�_�_o�_%o�/=o Oomoo�oo�o�o�o �o�o!3WE {i������ ���A�/�e�S�u� ���������я��� ��+�a�O���;o�� ��͟ߟ�o���%� K�9�o�����a����� ۯɯ�����#�Y� G�}�k�����ſ��տ �����C�1�g�U� w�yϋ��ϯ��ϛ��� �-�?�Q���u�c߅� �ߙ����������� ;�)�_�M�o�q��� ���������%��5� [�I��m��������� ������!E��] o���/�����/M�$T�BCSG_GRP� 2��  �M 
? ?�  x� t�����/��,/>+QX_d�@ �m!?M	 HBL>(M�&=$?B$  C�p�/��(}/�/Cz�/�-A��>(333?&f�f?��<%A��/@?0 >(�͘a6&5V0DHC?�=@��0=%1�5=$�1D"!!�?�?[?�?O�: �(&�(AETOO1OO��OgOyO�O�O�K�H�Q	V3.00~p	lr2d�C	*/P'TL>_�O3 aQ�I uPG]v_  �_�_�[QJ2X_Q�_�U�CFG ei l�Z�b��R�_Jh� Jopo~j"~o�o�o�o �o�o�o�o41 jU�y���� ���0��T�?�x� c�������ҏ����� �,�p� 7�I�[�� ��y���ğ���ӟ� ��0�B�T�f�!���u� �������M9	� ��-�c�Q���u��� ��Ͽ��߿��)�� M�;�q�_ρσϕ��� ��������7�%�G� m�[ߑ�ߵ��߇�� �ߛ��3�!�W�E�{� i����������� 	���S�A�w����� ��g��������� O=sa��� ����9' ]Kmo���� ���#//3/Y/� q/�/�/?/�/�/�/�/ �/??C?1?g?y?�? �?[?�?�?�?�?�?O -O?O�?OOuOcO�O�O �O�O�O�O�O�O_;_ )___M_�_q_�_�_�_ �_�_o�_%ooIo7o Yo[omo�o�o�o�o�o �o�/'�o�oiW �{������ �/��?�e�S���w� ����я㏝����+� �;�a�O���s����� ͟��ݟߟ�'��K� 9�o�]�������ɯ�� �ۯ���5�#�E�G� Y���	����˿u��� ��1��U�C�y�g� �ϯ����ϑ������ 	�+�Q�c�u�/�A߫� ���߽�������'� M�;�q�_����� ��������7�%�[� I��m����������� ����!3ݿK]� ������� ASe#5� �����//� =/+/M/O/a/�/�/�/ �/�/�/?�/?9?'? ]?K?�?o?�?�?�?�? �?�?�?#OOGO5OkO YO{O�O�O�O?q�O _�O�O_1_g_U_�_ y_�_�_�_�_�_	o�_ -oo=o?oQo�o�o�o �owo�o�o�o) 9;M�q��� ����%��I�7� m�[����������� ُ���3�!�W�i�_ ������O�՟ß��� 	���S�A�w����� ��k�ѯ��������  ?�C� �C�W�C��$TBJ�OP_GRP 2� �� _ ?�C�	o��v�"}�����@�� 0��  �� � � � �{C� @?����	 �BL  ~�Cр D]��������&�<��B$鰌���@��?�33C���X��f�q����'ϩϷ�;�2��G��@���?���z��_� �A5��ȍ�� �Ϡ����?�>�Q�4�F�;��pA��?�f�f@&ff?�ffWψ�� ��ߝ��P�������:v,�ƣ�?LQ�P�t�DH���� �@�333����>t�O�X�j�8���3Ꮁ���D"�������3�E��O�������9�� ���:�I�T�K���s� ]�k�������_��� ����)Z5��y�`}���C�C�C��ܱ��	V3.�0Ƴ	lr2d��*5��>�CN� E8� E�J� E\� E�n@ E��E��� E�� E��� E�� E�h� E�H E�0 E� E�e��� E�i�� E�x E�X� F�^D�  D�` E}_P Ee$mU0�;iGqR��^p Ekyu��r����(z�� E�}���X� 9�IR!�D%
M�3/E"C��I#��߄/k�ESTPARS 7����l�HR� ABLEW 1#}� C���(^' ��>)�'B�(�(B�J��'	�(E
�(�(�%C��(��(�(!�#RD	I�/���/�/�/??15�4O�?�;�?�?��?�?N�"S�?��  c:�O�O�O�O_ _2_ D_V_h_z_�_�_�_�_ �_�_�_
oob��@�O ���']iFOXOjO|O(?�:?L?^?p?�8�"CbN�UM  �*��ϰK�   ��"_CFG $�,{�c�@o�IMEBF_TT�!�e��� nvVER#oa�v�nsR 1%�+' 8@C�>��q �ho  ��� ��#�5�G�Y�k�}� ������ŏ׏���� V�1�C���g�y����� ����ӟ���	��-� ?�Q�c�u��������� ϯ���N�)�;��� _�q���������˿ݿ��"�q_&q�v@�u�� MI_CHAN�zw �u H�DBGLV��|u�u�!K��ETHERAD �?�%���I ��￷��ϓ(K�RO�UT�p!*J!������SNMAS�K�ȥs��255.Y�!W�i�{�!� �OOLOFS_D�I� �}�ORQCTRL &�{CJ/��T���/�A� S�e�w������� ������+�=�M����p�_����#PE_D�ETAIqȾ�PG�L_CONFIG� ,,y<q���/cell/$C�ID$/grp1��� 2DVC� �ρ�����j �#5GY�} �����fx/ /1/C/U/g/��/�/ �/�/�/�/t/	??-? ??Q?c?�/?�?�?�?�?�?�?gn}�?)O;O MO_OqO�O�a���O�M��?�O�O__(_:_ �?^_p_�_�_�_�_G_ �_�_ oo$o6oHo�_ lo~o�o�o�o�oUo�o �o 2D�ohz �����c�
� �.�@�R��v����� ����Џ_����*� <�N�`�������� ̟ޟm���&�8�J� \�럀�������ȯگ����User View ���}}1234567890�/�A�S��e�w��������2�|����� )�;Ϛ���
�3Ŀ�� �ϭϿ�����B�߲�4x�=�O�a�s߅ߗ��ϸ߲�5,�����@'�9�K��lﲾ6�� �����������^� ���7��Y�k�}������������8H��1CUg���� �lCamera����'BE�Qc u���������  �ù�9/K/ ]/o/�/�/:�/�/�/ &/�/?#?5?G?Y?���w��/�?�?�?�? �?�?�/#O5OGO�?kO }O�O�O�O�Ol?~7+� \O_#_5_G_Y_k_O �_�_�_�O�_�_�_o o1o�O~7+�_o�o �o�o�o�o�_�o! loEWi{��Fo ���4����1� C��og�y�������� ӏ���	��~7G��� U�g�y�������V�ӟ ���B��-�?�Q�c� u��~7�����ӯ� ��	��?�Q�c��� ��������ϿῈ���9m�"�4�F�X�j�|� #��ϲ���k�����ߠ�0�B�T���	�0 �Ϗߡ߳������ߐ� ��1���U�g�y�� ���V�h߮ �S�� �,�>�P�b�	���� ����������( ��+��t��� ��u��a: L^p��;uՈ; +��//(/:/� ^/p/�/��/�/�/�/ �/ ?���K�/L?^? p?�?�?�?M/�?�?�? 9?O$O6OHOZOlO? �`kO�O�O�O�O _ _�?6_H_Z_�O~_�_ �_�_�_�_O��{o_ $o6oHoZolo~o%_�o �o�oo�o�o 2<D�]  �Ys ��������x�'�9�   I Qo���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u��������=�  
�P(  ��gp( 	  ���߿��9�'�]� K�m�oρϷϥ�����t��źY� ̓o D�V�h��o�ߞ߰��� �����S3��"�4�{� X�j�|�������� ����A��0�B�T�f� x������������� ,>����t� ������� ]:L^���� ���# //$/k H/Z/l/~/�/�/�� �/�/�/C/ ?2?D?V? h?z?�/�?�?�?	?�? �?
OO.O@O�?dOvO �O�?�O�O�O�O�O_ MO_O<_N_`_�O�_�_ �_�_�_�_%_oo&o m_Jo\ono�o�o�o�_ �o�o�o3o"4F Xj�o�o��� ����0�B��f� x��������ҏ��� �O�,�>�P���t����������Ο���@ A����!�����۰��+frh:�\tpgl\ro�bots\lrm�200id[�_m�ate__�.xmlݟ��������ϯ�`���)����3� X�j�|�������Ŀֿ �����5�/�T�f� xϊϜϮ��������� ��1�+�P�b�t߆� �ߪ߼��������� -�'�L�^�p���� �������� ��)�#� H�Z�l�~��������� ������%�DV hz������ �
!@Rdv �������/t.:�p� ���E�<< C� ?�+[//S/u/�/ �/�/�/�/�/?�/? )?W?=?_?�?s?�?�?�?�?�?O��$T�PGL_OUTP�UT /#�#�/ ; CEXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_CE�; �@2345678901o-o?o Qocouo}c�o�o�o �o�o�o�o�o4FXj|z}��� �����,�>�P� b�t��������Ώ�� �����:�L�^�p� ���,���ʟܟ� � ��� �H�Z�l�~��� (���Ưد������ ��D�V�h�z�����6� ��Կ���
�ϴ�*� R�d�vψϚ�2�D��� ������*���8�`� r߄ߖߨ�@߶����� ��&��A}6!\�@n�������@=/�����C* ( 	  o2� �V�D�z� h��������������� 
@.dRt� ������@*`N�f�9  R&�����/� (/:/j�k/}//�/ �/�/�/�/�/Y/�/1? �/?g?y?S?�?�?? �?�??�?O-OOQO cO�?KO�O�OEO�O�O �O�O_uO�OM___�O g_�_o_�_�_�_;_o o�_�_Io#o5oo�o �_�o�oao�o�o�o 3E�o-{�'� ����W�/�A� �e�w�Q�c����� ������+���a� s�яw���C���ߟ� ˟�'����]���I� �����ɯۯ9�ï� #���G�Y�3�e���� ��ſ׿q�߿���� C�Uϳ�yϋ�%�w�����ϭ���	ߛ�$T�POFF_LIM� ��Мy���$�N_SV(��  ��:�P_�MON 0�)<�����2��$��STRTCHK �1�:�Y�B�VTCOMPATO����>�VWVAR �2o���S� ��� �3����$�_DEFPRO�G %��%?STYLE1+���_DISPLAY�/О�D�INST_�MSK  �� ���INUSER��߆�LCK���QUICKMEN��ކ�SCRE�����tpsc@����6�;�:�L�_P��ST��:�RACE_CFG 3o����3�	�
?����HNL 24S�x��� )��� %7I[m
��ITEM 25��� �%$1234567890��  =<��  !&��_����� ��>P/t4/ �D/j/���// (/�/L/�/?0?�/T? �/�/�/V? ?�?�?�? H?�?l?~?�?ObO�? �O�O�?�O O2O�OVO _zO:_L_�Ob_�O&_ �_
_�_._�_ oov_ o�_�_�_8o�_�o�o �o*o�oNo`oro�o �ohz�o�� 8�\�.��D�� ����������h� X�j�|������ďp� �����̟0�B�T�Ο x�$�J�\���h���� ���گ>����t�� ����s�ί��򯲿Ŀ (�ڿL���'ς�BϦ� R�xϊ���$�6� ��Z��,�>ߢ�b��� ����n߆� �����V� ��zߌ�U��p��ߔ�
��.�@�	���S��6����  �� ��e�\�
 r������=��UD1:\����� �R_GRP �17�� 	 @e�&F 4jX�|�� ���
������?�  ,>(^L �p����� / �$//H/6/l/Z/|/��/	��/�/�S�CB 28*� ?&?8?J?\?n?��?�?�?�UTOR?IAL 9*�����?�V_CONFIG :*���b����NO�=OUTPU�T ;*�?@��ZO�O�O�O�O�O �O
__._@_R_d_v_ <A�O�_�_�_�_�_�_ 
oo.o@oRodovo�_ �o�o�o�o�o�o *<N`r�o�� ������&�8� J�\�n��������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϓ��ϸ� ������ ��$�6�H� Z�l�~ߏϢߴ����� ����� �2�D�V�h� z��(O:E�O������  ��$�6�H�Z�l�~� ��������������  2DVhz�� ������
. @Rdv���� ���//*/</N/ `/r/�/�/�/��/�/ �/??&?8?J?\?n? �?�?�?�/�?�?�?�? O"O4OFOXOjO|O�O �O�O�?�O�O�O__ 0_B_T_f_x_�_�_�_ �O�_�_�_oo,o>o Poboto�o�o�o�_�o �o�o(:L^ p�����o��  ��$�6�H�Z�l�~�𐏢��������ӏ�ρ�����4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����+�>�P�b�t� ��������ο��� �'�:�L�^�pςϔ� �ϸ������� ��#� 6�H�Z�l�~ߐߢߴ� ��������� �1�D� V�h�z�������� ����
��-�@�R�d� v��������������� )�<N`r� ������ &7J\n��� �����/"/3 F/X/j/|/�/�/�/�/��/�/�/??-;�$�TX_SCREE�N 1<��π�}ip�nl/a0gen.htm-?�?�?�?�?��?%�Panel setup�<}��?OO1OCOUOgO�?�?�O�O�O�O �O�OoO_�O@_R_d_ v_�_�__#_�_�_�_ oo*o�_�_�_ro�o �o�o�o�oCo�ogo &8J\n�o�o� �����u�� F�X�j�|������ď ;������0�B����0>UALRM_M_SG ?M9�Z0 [�0*����؟˟ ��� ��%�C�I�z��m�����¯v�SEV7  ����t�ECFG >M5�W1  0%@�  A$�   ;B�0$
 ï7# M5W�i�{�������ÿ�տ����� �GR�P 2?
� 0�0&	 A�c�v�I�_BBL_NOT�E @
�T��l7"R09!��v�DEFPR�O��%�� (% ����9 �����(�� L�7�p�[߁ߦߑ��������l�FKEYD?ATA 1AM9M��p �0& �R�d��A���w�,(����0$����>��ANCEL�-����Q�8�EXT STEPZ�]��������ORE INFO ��������(L ^E�i������  �� � frh/gui�/whiteho?me.pngQ cu��(������//�FRH�/FCGTP/wzcancel< V/h/z/�/�/��/�/��/�/
??'/9#nextE/\?n?�?�?�? �/�?�?�?�?O"O-?7#infoK?bOtO �O�O�O�?�O�O�O_ _(_�OL_^_p_�_�_ �_�_G_�_�_ oo$o 6o�_Zolo~o�o�o�o Co�o�o�o 2D �ohz����Q ��
��.�@�O� v���������Џ�� ��*�<�N�ݏr��� ������̟[�ޟ�� &�8�J�\�럀����� ��ȯگi����"�4� F�X��j�������Ŀ ֿ�w���0�B�T� f����ϜϮ������� s����,�>�P�b�t� ߘߪ߼������߁� �(�:�L�^�p��߂� ��������� ���$�@6�H�Z�l�~�U�����$����������������, �=�aH��~ ������9 K2oV���� ���/#/
/G/./ k/}/\��/�/�/�/�/ �/
�?1?C?U?g?y? �??�?�?�?�?�?	O �?-O?OQOcOuO�OO �O�O�O�O�O__�O ;_M___q_�_�_$_�_ �_�_�_oo�_7oIo [omoo�o�o2o�o�o �o�o!�oEWi {��.���� ��/��S�e�w��� ����<�я����� +���O�a�s������� ���/ߟ���'�9� @�]�o���������ɯ X�����#�5�G�֯ k�}�������ſT�� ����1�C�U��y� �ϝϯ�����b���	� �-�?�Q���u߇ߙ� �߽�����p���)� ;�M�_��߃���� ����l���%�7�I� [�m������������ ��z�!3EWi ����������А��А���$6H j|V,h/�`/�� �/�+//O/a/H/ �/l/�/�/�/�/�/? ?�/9? ?]?D?�?�? z?�?�?�?�?̟O#O 5OGOYOkOz�O�O�O �O�O�O�O�O_1_C_ U_g_y__�_�_�_�_ �_�_�_o-o?oQoco uo�oo�o�o�o�o�o �o);M_q� ������� �7�I�[�m���� � ��Ǐُ������3� E�W�i�{�����.�ß ՟�������A�S� e�w�����*���ѯ� ����+�OO�a�s� ��������Ϳ߿�� �'�9�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� ��T�������1�C� ��g�y������P� ����	��-�?�Q��� u�����������^��� );M��q� �����l %7I[��� ���h�/!/3/�E/W/i/@�k+�>@�����/�/ �-�/�/�/�&,�?? �?A?(?e?w?^?�?�? �?�?�?�?�?O+OO OO6OsO�OlO�O�O�O �O�O_�O'__K_]_ <��_�_�_�_�_�_� �_o#o5oGoYoko�_ �o�o�o�o�o�oxo 1CUg�o�� �������-� ?�Q�c�u�������� Ϗ�󏂏�)�;�M� _�q��������˟ݟ ����%�7�I�[�m� ������ǯٯ��� ���3�E�W�i�{��� ���ÿտ���Ϛ� /�A�S�e�wωϛ�r_ ���������� �=� O�a�s߅ߗߩ�8��� ������'��K�]� o����4������� ���#�5���Y�k�}� ������B������� 1��Ugy�� ��P��	- ?�cu���� L��//)/;/M/ �q/�/�/�/�/�/Z/ �/??%?7?I?�/m?�?�?�?�?�?�?����;������OO(M OJO\O6F,H_�O@_�O�O�O�O �O_�O/_A_(_e_L_ �_�_�_�_�_�_�_�_ o o=o$oaosoZo�o ~o�o�o���o' 9KZ?o���� ��j��#�5�G� Y��}�������ŏ׏ f�����1�C�U�g� ����������ӟ�t� 	��-�?�Q�c�򟇯 ������ϯ�󯂯� )�;�M�_�q� ����� ��˿ݿ�~��%�7� I�[�m��ϣϵ��� �����ό�!�3�E�W� i�{�
ߟ߱������� ����o/�A�S�e�w� ��߭��������� ���=�O�a�s����� &����������� 9K]o���4 ����#�G Yk}��0�� ��//1/�U/g/ y/�/�/�/>/�/�/�/ 	??-?�/Q?c?u?�? �?�?�?L?�?�?OO )O;O�?_OqO�O�O�O �OHO�O�O__%_7_�I_ �K[� ����t_�_�]p_�_�_�V,�o�_�o!o oEoWo>o{obo�o�o �o�o�o�o�o/ SeL�p��� ����+�=��a� s����������Oߏ� ��'�9�K�ڏo��� ������ɟX����� #�5�G�֟k�}����� ��ůׯf�����1� C�U��y��������� ӿb���	��-�?�Q� c��ϙϫϽ����� p���)�;�M�_��� �ߕߧ߹�������~� �%�7�I�[�m��ߑ� ���������z��!� 3�E�W�i�{�R����� �������� �/A Sew���� ���+=Oa s������ //�9/K/]/o/�/ �/"/�/�/�/�/�/? �/5?G?Y?k?}?�?�? 0?�?�?�?�?OO�? COUOgOyO�O�O,O�O �O�O�O	__-_�OQ_ c_u_�_�_�_:_�_�_ �_oo)o�_Mo_oqo��o�o�o�o���k}�������o@�o}�o*<v,(� m ��x���� ��!��E�,�i�{� b�����ÏՏ������ ��A�S�:�w�^��� ����џ�����+� :oO�a�s��������� J�߯���'�9�ȯ ]�o���������F�ۿ ����#�5�G�ֿk� }Ϗϡϳ���T����� ��1�C���g�yߋ� �߯�����b���	�� -�?�Q���u���� ����^�����)�;� M�_������������ ��l�%7I[ �������� !3EWip �������� ///A/S/e/w//�/ �/�/�/�/�/�/?+? =?O?a?s?�??�?�? �?�?�?O�?'O9OKO ]OoO�OO�O�O�O�O �O�O_�O5_G_Y_k_ }_�__�_�_�_�_�_ o�_1oCoUogoyo�o �o,o�o�o�o�o	 �o?Qcu��( ������)� �+�� ���T�f�x�P�������,��ݏ����%� 7��[�B����x��� ��ٟ�ҟ���3�E� ,�i�P���t���ï�� �ί���A�S�e� w��������ѿ��� ��+Ϻ�O�a�sυ� �ϩ�8��������� '߶�K�]�o߁ߓߥ� ��F��������#�5� ��Y�k�}����B� ��������1�C��� g�y���������P��� ��	-?��cu �����^� );M�q�� ���Z�//%/ 7/I/[/2�/�/�/�/ �/�/��/?!?3?E? W?i?�/�?�?�?�?�? �?v?OO/OAOSOeO �?�O�O�O�O�O�O�O �O_+_=_O_a_s__ �_�_�_�_�_�_�_o 'o9oKo]ooo�oo�o �o�o�o�o�o�o#5 GYk}��� �����1�C�U� g�y��������ӏ� ��	���-�?�Q�c�u�h����p ���p ���ğ֟���
����,�M� � q�X�������˯��� ��%��I�[�B�� f�������ٿ����� !�3��W�>�{ύ�l/ ������������/� A�S�e�w߉ߛ�*߿� ���������=�O� a�s���&������ ����'���K�]�o� ������4��������� #��GYk}� ��B��� 1�Ugy��� >���	//-/?/ �c/u/�/�/�/�/L/ �/�/??)?;?�/_? q?�?�?�?�?�?���? OO%O7OIOP?mOO �O�O�O�O�OhO�O_ !_3_E_W_�O{_�_�_ �_�_�_d_�_oo/o AoSoeo�_�o�o�o�o �o�oro+=O a�o������ ���'�9�K�]�o� �������ɏۏ�|� �#�5�G�Y�k�}�� ����şן������ 1�C�U�g�y���������ӯ���	��$U�I_INUSER  ���*���  �
��_MENH�IST 1B*��  (� 7���(/S�OFTPART/�GENLINK?�current=�menupage?,153,1I���8ο��� ����962��>�P�b�t���'�36-����� ���χϙϫ�@�R�d� v�ؓߥ߷������� �ߎ�#�5�G�Y�k�}� ������������ �1�C�U�g�y�������~���������� �9K]o� �"����� ��GYk}�� 0����//� C/U/g/y/�/�/,/>/ �/�/�/	??-?�/Q? c?u?�?�?�?�����? �?OO)O;O>?_OqO �O�O�O�OHO�O�O_ _%_7_I_�Om__�_ �_�_�_V_�_�_o!o 3oEo�_io{o�o�o�o �o�odo�o/A S�ow����� �?�?��+�=�O�a� d��������͏ߏn� ��'�9�K�]�o��� ������ɟ۟�|�� #�5�G�Y�k������� ��ůׯ������1� C�U�g�y�������� ӿ�����-�?�Q� c�uχϊ��Ͻ����� ��ߔϦ�;�M�_�q� �ߕ�$߹�������� ��7�I�[�m���  �2����������!� ��E�W�i�{�����.��������������$UI_PAN�EDATA 1D����S�  	�} � FRH/FCG�TP/FLEXU�IF.HTM?connid=0/������)  grim��  d  $6HZl�~ ������� / /D/V/=/z/a/�/�/��/�/�� � �"	? ?2?D?V?h? �/�?��?�?�?�?�? 
OO�?@O'OdOKOvO �O�O�O�O�O�O�O_@�O<_N_5_r_�,�V U�?�_�_�_�_�_o b_3o�?Woio{o�o�o �oo�o�o�o�o/ A(eL�p�� ������_�_O� a�s��������͏@o ���'�9�K�]�ď ��h�����ɟ۟�� �#�5��Y�@�}��� v���&�8������ 1�C���g�y�쏝��� ��ӿ���^���?� Q�8�u�\ϙϫϒ��� �������)��M��� ү���ߧ߹������� B�7�I�[�m�� ���ߵ��������� !��E�,�i�P����� ����������l�~�/ ASew���� � ���+=� aH�l���� �//�9/ /]/o/ V/�/�/�/�/�/ ?#?v/G?Y?�}?�? �?�?�?�?>?�?�?O 1OOUO<OyO�OrO�O �O�O�O�O	_�O-_�/�/}�>_w_�_�_�_�_�_)e_�_i5�_"o 4oFoXojo|o�_�o�o �o�o�o�o�oB T;x_�����b8�#�+�$UI_�POSTYPE � �%�� 	 �5��Q�UICKMEN � �"�8��R�ESTORE 1�E�%  O��k2������k2mڏ��'� 9�K��o��������� Z�۟����#�Ώ0� B�T�Ɵ������ůׯ z�����1�C�U��� y���������l�ο� �d�-�?�Q�c�u�� �ϫϽ����τ��� )�;�M����l�~��� �����������7� I�[�m��"����� �������
����W� i�{�����B������� ����ASew��C�SCRES�?�X�u1s]c��u2�3�U4�5�6�7��8��TAT��� g��%�zUSE1R� ��ks�WU3W4W5W6W�7W8W�NDO_CFG F��NPMQ�OP_CRM5  IU���PDA��NoneF�8_INFO 1G�%5	 e�0%�$/ b8/S/6/w/�/l/�/ �/�/�/�/??�/=?�O?2?s?<��OFF?SET J�!�?*��2�?�?�? �?'OO0O]OTOfO�? jO�O�O�O�O�O�O#_ _,_>_�Kh��]x_�_�
�_�_�8UFRA�ME��SRTO?L_ABRT�_��bENBohGR�P 1K��d�Cz  A�mcka,@ko}o�o�o�o�f�o��ojR�U7h�&kMSK  :e	!&kmN�Q%)�%Z_�{E�VARS_C�ONFI�L�; �FP*��xCM�RSb2R�;�y, 	��p`01�: SC130E�F2 *�
�*��OX��t�� V�?��`@�`p�`��~ �_^� h�#����ȏ�qÏ��Za��eA�,܏�-�, B���H�,L�ԏm����� `�����ٟğ����� 3����i�T�f���R��ïկ�tISIONOTMOU`:t���쥙SS��S�0ba� FR:\�\��A\گ ��� UD1-�LO�G:�  S�EX�_�,' B@ ����r�j���r�ÿ�* �� n6  ��q�#��t�`�����  =����5�*2�s�TRAI�N����D¿P  d�y�p5�"���rT�=(��5Ž�V����� ������4�"�8�F�X߀j�|ߎߠ���W��_��RE�UZi�r�t/LEXE�V�|��1-��~MPHA%S	��D��s�RTD_FILT�ER 2W�; �RU�U�������� ����&�8�J��J�� {�����������������vSHIFT�r1X�;
 < ��iwV|�� ����!�
0 i@R�v����	LIVE/S�NA�s%vsf�liv;����� �0U�p
"menu /%/��/�/m"�6�YE	Gr2MO��Z'���`�$W�AITDINEND��#x�$O7p7���*?S>?9TIM.8u��i<G�/�= ?�;=?�:\?�:{?8RELER�8o�$��<��!_ACT�=H8CxrB6� [\{�/x�O�VrBRDIS�p�9o�$XVR��\'��$ZABC�Sc]� ,�X2��O�]ZIP�^�����_�_�_TZM�PCF_G 1_Zk 0s�~_o�W�Sc`Zi@q�� �8��Ro�a<+�Wo �o�oAo�oeiH����o �o�o�o�oA�ot�D��I����� ��{P�P�aj_S�bPYLINDx�b��[ � �,(  *\�m���Y���}����� o���� V�7���[�B�T���ԏ ��ǟٟ�����~�3� �W�>�������S[ cs2c�W�A ��_ ����n#��G�Kyhگw�Kw���A�*��SPHERE 2d<���ͿA�ƿ� �'�o���]�o�럓� 2���ϰ�����F�#� 5�|ώ�k��Ϗ�v߈����������PZZ\F �HF