��   �A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����BIN_C�FG_T   �X 	$ENTR�IES  $�Q0FP?NG1�F1O2F2OP�z ?CNETG����DHCP_C�TRL.  0{ 7 ABLE? �$IPUS�R�ETRAT�$SETHOST��NSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!� FT� =@� LOG_8	,�CMO>$DN�LD_FILTE�R�SUBDIR'CAPC����8 .. 4� H{ADDRTYP�=H NGTH��f��z +LSq� D $RO�BOTIG �PE�ER�� MASKn�MRU~OMG�DEV������PINFO� � $$$T�I ��RC�M+T A�$( /�QSIZ�!S� TATU�S_%$MAIL�SERV $P�LAN� <$L�IN<$CLU���<$TO�P7$CC�&FR�&Y�JEC|!Z%EN�B � ALAR:!B�TP,�#,�V8 S��$VA5R�)M�ON�&����&APPL�&PAp� �%��'POR��Y#_�!�"ALER�T�&i2URL �}Z3ATTAC���0ERR_THROU3US�9H!�8�� CH- c%�4MA�X?WS_|1���1MOD��1I��  �1o (�1PoWD  � LA��0�ND�1TRYFDELA-C�0G'AERSI��1Q'�ROBICLK_HM8 0Q'� XML+ 3_SGFRMU3T� f!OUU3 G_�-COP1�F33�AQ'qC[2�%�B_AU�� 9 R�!UPD�b&PCOU{!�CF�O 2 
$�V*W�@c%ACC�_HYQSNA�UM�MY1oW2"$DM�* $DISL��SN,#	3 ��	o!�"%"_W�I�CTZ_IND9E�3�POFF� ~UR�YD��S�  
 t Z!KRT�0N�(cD�.)bHOUU#E%A/f�Va>fVaMfLOCAܗ #$NS0H_[HE���@I��/  d�PARP�H&�_IPF�W�_* O�F�PQF�AsD90�VHO_�� 5R42PS�a?�wTEL� P����90WORjAXQE� LV�O#�FS1�ICEد[p� �$�c  � zq��
��
�op�PS�Axw�# �i�qIz0A�Lw�q'0 �x
�
��F�����p�r�uw�$� 2�{���r#���� ��}��!�qi����$�� _FLTR  \�y�p ���������}�$�}2�}��bSHAR� 1�y Pe���t
�G�6�k�.���R� ��v�������П1� ��U��y�<���`�r� ӯ�������ޯ?�� �u�8���\������ ��ڿ��;���_�"� ��FϏ�jϸ��Ϡ�� ��%���I��m�0�B� ��f��ߊ��߮���� ��E��i�,��P�� t���������/����z _LUA1��x/!1.j�08����i�1z���2551.��q�����uh�2o��������������3����^ 1C��4_��� ������5���N�!3��6O��� u������QJ������ �(�?� Q� '��<a/�/�/{/�/�/�/�/?&?��P?V?h? z?9?�?�?�?�?�?�?
OO��?���ufO�QL
ZDT Status�?uO�O��O�O��}iRC�onnect: �irc�D//alert�N&_8_J_\_ �G�O�_�_�_�_�_�_����sP 2ـd���_o1oCoUogoyo �o�o�o�o�o�o�o�s�$$c962b3�7a-1ac0-�eb2a-f1c�7-8c6eb5�f01a8c  (y_J�On���R���ـP(�X" �rZJ�u3 �v[C] )�,$e"�ـ[��M� 4�q�X�~�����ˏ�� ���%��I�0�B���f��������w��W�8 DM_=!yW�G�SNTP咋	�%��-���>������K�4#���USTOM �
�F��W  |�3$TCPIP撅�XHO%S"��E�LO�W�T!�E�H�!Tb���rj3_tpdQO� \��!KC�L�������v!CRTY�G���O"(�!CONS��� ��ib_smon����