��  	NK�A��*SYST�EM*��V9.1�035 7/1�9/2017 �A  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  ����AIO_CN�V� l� RA�C�LO�MOD�_TYP@FIR��HAL�>#INw_OU�FAC� �gINTERCEmPfBI�IZ@�!LRM_REC�O"  � AL]M�"ENB���&sON�!� MDG/� 0 $DEBUG1A�"d�$�3AO� ."��!_�IF� P �$ENABL@�C#� P dC#U5K��!MA�B �"�
f� OG�f d �PPINFOEQ�/ �L A q?1R5/ H0�f69EQUIP� 20NAM�� ��2_OVR��$VERSI�� �!PCOUP�LE,   $�!PP_D0CES�0�!�81�!"PC�> [1	 � �$SOFT�T_�ID�2TOTAL7_EQ� $@%@�NO(BU SPI_OINDE]=EX�2SCREEN_�4��2SIG�0��?�;@PK_FI�0	$THK�Y�GPANE0D �� DUMMY1"d�D�!�E4�A!�RG1R�
 � _$TIT1d  ��� �Dd�D� �D�@��D5�F6�F7�F8
�F9�G0�GW�A�EW�A�E.W18W �F�LW1VW2aR!SB�N_CF�! 	8� !J� ; 
2f1�_CMNT�$�FLAGS]�C�HE"� � ELL�SETUP �� $HO�0 P�R<0%3cMAC{RO?bREPRHhD0D+<@�bb{jd^ UTOB U��0 9DoEVIC�CTI�0��� @13��`B�ce#VAL�#IS�P_UNI��`_�DO�f7�iFR_FZ@K%D13�A�c�C_WA�d�a+z�OFF_�0N�DELXxLF0�a�Acq��b?�adp�C?�1`yA�E�C#�s�A�TBXt���MO<� XsE � [�MXs���qREV��BIL�w19��AXI� �rR 7 � OD5`��$NO�PM@��p�
� �/�"`�� +�V�  ��X@D�T p �E RD_E
��q�$FSSB�&$CHKBD_SE�e�AG� Gj2 "_��TB��� Vxt:5p}�C �a_EDu >� � C2�eA`S8p�4%$l �tt$OP\@B�bq!�_OK��US�1P_C� !��d��U S`LACI�!�Rae���� �aCOM9M� �0$Da�w��H@dp ��O�B�IG�ALLOW� �(KD2�2e@VA�Rݕd!PAB =m��BL#@S � ,�K�a��`S+p"@M�_O]"���C�CGXpN�!o $��_ID�L�`��$�� B��)AS� c�CCBD	D�!{�I����LPz�|84_ CCSCH�1�` OOL��`�M�M��S�C�s$MEA�P\t�`Tg`�!���TRQ�a�CN����FS3k��!/0_F��( )��p���U� �!B �CFn�T X0GR�0���M�qNFLIx�u�@UIRE�x���!� SWIT=$�(�N'`S�"CF_��G� �A0WOARNM pP���r�PLX��NST� �COR-���`FL{TRܵTRAT �TR�� $ACC�a�� �r$OcRI�.&��RTj`�_SFg CHG*x@I��Tp�A
�IF�T�!���>� � �#a����HDh�Rq��2B�BJ; �C����3��U4��5��6��7��e8��9�!h�CO�S <� i�{���x3�2-�LLEC��}�rMULTIr�
2ʓyA
2FS��I�LD	�
1v�B@T_��R  4� S�TY2pbܖ=�)�2ܐ��`��0� |A06$��`@�ޔa`�* ��TOx�:�E,�EXTB�e�p?��Be�f22n0,����0��R�.'�������� �"�/%9a9�����cg����� ���A�C�?�ME� �� q�Ջ��! L0���� ��cpA��$JOB�Ȱ�l�K�;IG��" d{�^� p�����-'��8�嗷��ACO_M��b#� t{�F� �CNG�AiBA� w�DɁ M
/1Bk�j0W�F@�yP�`zm÷$ϰ$��t�a�"��
2J"�_R�a"C��J%���J�D/5CԽ��Fn@b �W�P�O�л!% \0RO�6i(��S��O_NOM_ �`n#�jc�Aᦰ������ T0�&"�@<�U��Pk��e�RA@@n �3"��?�
$TF�<�D%3S�TP�pU�1���%�%�H�b�T1Y*E������#��p�%���A�YNT�"�TDBGDE�!'���PU�@��=�82C�AX�㟲[uwTAI�cBUF��8+ѳ!\1( ����&��PIӄ'�P�D7MC8MP9� S6F>D7SIMQS�@�wKEE�3PAT ���"�"#�"m�A�Cb%)���pw`JB��U�vaDEC�:[�58*�A�$* �����v�MP��$G- �G��_e jc��1_�FP�e TCJFS W�MEb��_D?#� J��V��V��Q��FJR�F�V�SEGFRA�6�O����@T_LsIN���CPVF�q;��`t �$+G�l��B�����B"r�2�,` +,��ܵQ�� F�P�0'`�bRTm�aY�1SIZ��r�}T\V�TgS- �Z�YQRSINF� ІC�@�@�I�\�@�Xk@�@Le�8d )@fCRC��?sCC�e�@6hJA�� JBۢqdeJA�Hh�Q"eD����|iC�kcp���~D�`���f< �hE�V�f�F�a_}EFo@Nv�@�1ܶ�h+�,݀�C%�+d!V'SCA��e Ajv��Rɰ1�C�-��	��MARGh�C&�F�@6�_AD�Q��_@LI����kb`���8J|��#`r�.� <�Nߌ�S�t5��� �HANCq�$LG��O���{�4 ��B(�A�< ��0R�rrC~�ME�1���)0fy�RA��~�AZ��ň�`@%Oa�FCT h��p)���eb_@�0� ADI�O���A ��<X������L�S���B�BMP��D�PY�7A4�AE�S�P�cB H�U�0M�MENU�/��T#IT�q���%��AH�!)1��L�Ѐ�0d,�Q��OR	R$����	P  ��Ou���O��4%�������E�V/#(У DBPX�WO�P��1)�$sSK�2itp��T9�TRL�2 ��� AC�@A�&�I�ND� DJ8��_�kp1��;���PL�	Q�2WA��ΠE"(�D�!ۧ�!�R�>��UMMY9"��m1�� �DBρ��3c�)1PR�Q� 
�������4 ���'$��$^�Q �L<�5I��[�c���6o�����PC�7����EN�E��q8�����RECOR��9�H&�C#� 74$L��5$<�2�����@���A�_DJ�?0ROS� 2�À{�mӽIñ�;�a�P�A/��BETURYN_�gcMR��U� v��CR.�EWM�B=�0GNAL� 2�$LA]�Ş6{$P��7$P�F��8���!M`C�����DO�@��)��|Kb/�GO_AW���@�MOޑ:��� ��DCSS_CN
��Y��:Y��T@���Z�ID'��2]�2
k�N�O��D��`�I:� ; P �$��RBoR�P�Ik�PO��I_B�Y!�����T�RD�H�NDG��< <��A��c@�SO DSBL��S�6�l���F�;LS�q= H��0<60k�TOFBm�$FE9����l�Dө�q>b�DO7A,S`�MC@��[��4���ʚ�H�W( �MY�7��SLAV�r?�BIN� ��63�֭�_�@P!P�`@ ���А��А�u��!"��Z�?�Y�I$�����W���NTV�3[�VE4�SKAI��A��3��2�B�7AJv7A��~DSAqF�ZE_SV.��EXCLU�� N�rONL��>Y���]��EA�HI_V�I���PPLYӠRb�sH\0Q�l_M$"}��VRFY_��zjM�s$IO�0���#`1�B���O���oLSp����4��!�l��@�P�K�$J��AUTOCN� ��4l���N[WCHD\�5�_�l���AF9�CP��TT�!�=�6�j� #AӰf�\!_@w g ��;�SGp� B �* CUR����1� �� �@��F��F��ANNUN��=#l�������d�1).!#`6*�R&�EF�I��C� @�F"Ŕ`OT����������n M��NIC�D�T��",W� AU��$D{AY�LOAD�����"�5�#EFF�_AXI\�EӰęQ��O0����_RwTRQ�qF DWq�H0�RT3@\45 2E�@�wC1��� �A�p81�qG 	0K!�1A�T�2�/��DU��/��|�CAB�qH|"�p@�0P@ID�@PW�s�5@Q_@V��V_�0z0Ҁ��DIAG��qI?� /$V��YUT�GHA�Q��NJ��R�Rʲ�!�TVE� SW�A���P�0��BC5z0F�PC1OH�Y5�1PP�@ cIR���RB�P�2�3�q��8 aL �BBAS;�G@��Ҁ�E���5z0H�xH0J��URQDW�EMS�@HUAKp�EsB�TLIFEkpT#rP�~RN�Qb�U.!�S�bZq��."C���3�N��Y�p��FL�Ah�/ OVJ��VH�E��BSUPPO$����~R��_�T���Q_Xw�d.�)gZ&jW&j��)g�.!'��.�XZ��3��QY2��hC �TF�G�MEN��pKD.pn)@CT�?�J `��CA�CHE%w�bSIZдV�PH��N��UFFI%`Z�kt��2�6�S�MSW�eK 8�KEYoIMAG��TM!����Kq��Fv�8�O�CVIE�@�L �� �L���w�?�� 	 C�6��M�P0��ST��! �r堻t�t0�t0>�pEMAILp�\�x�!�qFAUL�"qN�rZÖ�COU��䃐9�T�2AO<' $&���S�0�0;IT��BUF�gw�P�g��Ӑɐ�PBR����Cv�A�'���4�SAV��_�d@�bw�F���'�2&P�����D�5�_R���� ��OTN�V�3P� ����( �n�h�F� XR�C�у_G�S
�YN)_�A5pP�2D�ճ�����BM�2�PT
�F��0��(���4qQ�` Gs��!&��+��������4qR�������C_E���KU��� ���RCq����DSPl[v�PCF�IM�� =�c�x�<@U��PTř �pIP����A7D  <�TH렋��0�#0TH�=�HSD=I:�ABSC���`ɰVM����#��34NV*G��`$:�R�F�Aj�d����G���SC.B����M�ERe�FBCM�Pe�ET� mS9rFU`DUF�0p��vb0CD3���l����o�NO4
4qTP0��޲�%ܴV�%PS۵C���	C7!�1ٳ'�5p_UH *�LR� ���&�h�P W��^� �\Ʈ!\�1\�1\�T#q\�7Y�8Y�9Yʨ�P[�e�1r�1�1���1��1��1��1*��1��2��2e�r�U2�2��2��2��U2��2��2��3�ʥ3e�3r��3��3���3��3��3��32��4��XT?A4qV <�������V���VŌ��� �'@FD�R.DWT2�V��~R���~RRE�Mg@Fq��BOVM���A�TROVf�DT��4�MXC��IN��P3�+AIN�DR��R
~�ޠj�$DGR��C=�p�UrtADX6=�RIV���R�BGEAR�I%OkEK�TN�����1iXa gp`�SZ_�MCMy`~Q�Fv�PUR��X ,鱞u�? �Pz?�P �A?PE@� X�1��t���Y0j3PP:�;@RIµ��p_�ETUP2_� Z 0^�TD �����h��"��_�BACv�[ T(�p_�ɔ)Ú%�#!����IFI�A��t��E��@PT�Bl�F�LUI�d\ � ��w(�UR Q���R@����U�CCh0I��u$�S@?x��JƐCO��VR�T��� x$SHO8g1= �ASSΠ�8�U����BG_�� ��������´�^IDATA2A]�KFU;1��5$2��p��J�`2A^ |��wNAV*���ʼ� �S�r�S$�VISI��SCF*�SEv ��5V� O�1/1B'e=@^�&$PO� I�A�FMR2��_ ��Ͱ�2 ��א�&����+�(��U�_����h@GIT_:��f@M��|����DGCLF�EoDGDY�8LDhB��5�V���T !M���s`!�O9 T��FS���ta P��+Bדj�$EX_+ABH+A1F�9��Rj,@3dK5dF�G���%b �` ��SW���O9VDEBUG���A	�GR� �Un[�BKUf�O1.�7 �0PO30�I��@���E�@M�LOYO:�QSM_0E���!p�P_E c� x@���ATER�M4Ud=U!ORI䷑9Pe=U��SM_�Đ�9Pf=U����* |XgVV5 UP>}rh� -o�2�c�KS�Pd� G��Z�0ELTO�q�$USEs�NFIG�b�Q; �A��bT�T�e$UFRʒ�$߰�Q&`��j0OT�3g"�TA͠��EcN;ST��PAT¡�`�[bPTHJ��Ep�pԂ���RARTŀ��U�Ł�r�QREL<�ja�SHFT���Qaa�h_�R����zV% �P$�W�`g�1��8�x�a�SHI�`�4�U� ��AYLO ��Z�p�My �aaV!󵿠ERVd�,q� �h��Ag���b�,�u��,RCx�AScYM����QWJg���E��a�y���U�t��p��e�0{v�eaPv�Ip&�vOR���M�#��@#Q�$i�1"�B	V`` `Y�� H9O�Dj �Gb0,� ͰOC�Q�A!$OP�$F�J�F� ��� �2��R:�a�OU�acerR_e�Ɉ�a��e$PWR��IM�]rR_���d� {Ptc�QUD�  y����k� $Hȕ!^n�ADDR��H&QAGcb��|�u�-�R�".Al H��Sa��!�㴕㴕ô���S1ES1�#� HS���#�m $3 ��_D����@���PRM_�f"!HTTP_�ްHAn (�OcBJ� u��$���LERcw�1�� o � �痡AB_�TS��Sm��\�KRL$�HITCOU�����!ƀ������ƀ.ǀSS���W�JQUERYO_FLA�Qw�W����QAp���IN'CPUxB�!O2����d�I�ʔJ�ؔJ���_�IOLN�q���k0C�!$SL��"$INPUTM_)Q$䀙�P�#w Cu�SLA�1 r����ѵʹ��s���r!IO�F�_ASBs� $ALW��aN�UzP��`ae���@��.pH�Y��P�)�EQ�UOPEt `�n���@b�@�b�GƘ���P�� 䀎ǲ�Gƿ¨ƫQ� 9M�qRu l\@s�TADr^�A�TI����:�30ի`PS6�BU30IDW0�� �7�Ԁ6�p��2�S`vȲ��#����N��30���IRC�A���� w �� ��1�Y��EA 8��џ!��b��ׇ�R{`�q9��DAYy_?�:�NTVAa�N�&���e2�&�SCA>p&�CL��?���?Ҝ RxjߋԀb,�ա�N_��C2��?��SyȲ( ���ဦ�R�?�6���(! �2x� ���Rzp��R��LABSa�+�301�UNI4�ePITY������UJR�%{ ����FU@
w�g��D^s�$J7��O�r/$J8��7d@�$����70���8����oAPHI� Q��z��D-@J7J8�� L_KE\� o �KK�LM��� | <ʰXR��?��WATCH�_� Fs��ELDb	y� 3E} f0�IaVRp�֓CTR`�c���B� LGO�~� !��LG�Zw�@�@���FD�I��Q ��6P�� ��� @����6P�p�p�E�P�!_CM7c�T@�A1F�q���� �(��b ��@���'I�(P�6P�� �RSV p`  (�s�LN���"z�����@TAҲ" t!��U���!m�L�#�"DAU�%EA �4 ���"Ƴ GH��.Q�BO�O���� C/�4�IT��$�0+�sRE��8SCR�,��0�DI*�S `�0RGI)R�0=;��#Ð��f2¤�Sc��WpD4��$#�JGM�7�MNCH��FNt)�6K�7PRG�9�UF�8p�8FWDv�8HLISTP�:�V�8eP�8� �8RS"@IH#��; �CtC �r#�Q�x7�IU��4@w7��5� 8��2G�9�`PO�G#J35C��4OCU�HRGE]X�TUI�5I< ����<�dQQ�3[S�0\��`?��	[�%5�`v$1NOTVANA��R=�AI1�|�l�uDCS༓�Sʓ�RO�XO�WS��b�X9S h[8IGN� ?���1����TDEVzGLL�qm!c L���i�� m�T�$��d�:��W�CAd��� ����E�'��*�@1�e2�e3�a��8R�P��� ����b�T��5��7�Q����@6��;vST��R� Y6��P^p �$ElvCl{����{v�vw�T��� L ,�>���S�5�SǶ����8�EN �8��#"5_ �	�i�%�X�%0��MCu"�� ���CLDP|���UTRQLIU�p�S��Q�?�FLGgr?� �s�j�D�s���LDs�]�s�ORG0��vB���RE0����҄ʓ҄ؒ 0� �� � 	\�wEN�s�SVe Q�, �����,�4�RCLMC�B�ҏ�T�o�4�� M袠�� �@ $DEBUG���R��T�P-�E��Tgq���ISCv�� d�~!qRQ, 	�DgSTBO0F� ��D1	�AX�R. �%�_EXCES���RߒM���������Tl!ߒSCp �*��� �_�����Б�#�5���K�� �\,���O0��B�L�IC�tB0QUI[RE�CMO�O�����p���L�pM�� �0�<��ݣR��� MND�!� C�|"s"�{�D�>�$INAUT51�$GRSM��,`Ngr�o�Ca���g�PS�TL�� 4��L�OCvRI>@uE�X��ANG�R���[��oAQ���1-��MF� B�8y�r�@�uh�p ��gSUP�uW�FX���IGG1 � ���soV��r�F�tb  %\s��_p��_p �ư��C�g������`I��� Mt0�MD-�K�);��PF�Y�C�H���F��DIU�F�ANSW�j1FԵa,QF�D�#)�e�Ou�*�� � d�CU� V��u����.�O]1_���� ����s:Ö�/�����P��K@#p��P���KE�B_ �-$qB����pND2[G�2_TX�tXGTRA�Ss�m��<�LO� � �b�����	��y�ҩ��ے�RR2v��0 �#��!A1� d�$CALI2�pGt�Q��2�`RIN����<$R��SW0�`�#�m�ABCA�D�_JY�����:�_Ju3N�
H�1SP� $����PH�o�3n����p����Jm����)�OvaIMm�4�CSKP`�������	J�!4�Q�����_AZ0���@�EL[a���OCMaP�5�Pq� RTʑ�k��1�����2p1і�|P�
Z�SM�GZ@�2�JG�S�CLE��SPH_@`4���_������RTER"�����INACp�����^2����p_N���8=q4�̠45}��BDIV��Fm DHE�u����`�$V�����|Q�$� �́�`�_��ذR�ӡ��H �$BELQ ����_ACCEL�Q��m��IRC_R4�n�ŀNTPq<sO$PS�D�L� N $$Y�'�!�P@&>��['�['3*"��H�_�a�� �!/�r�C? �_MGoQ�$DD�! 42$FW����%����(DE�+PPA�BN2'RO� EE �"�a?Q��a������� $USE_����SP��C�@�SYh0�/� �qYN�AA�y6��]�y1M������R� OLK#�4INC����"�$	��7<��
�ENCS���`��"!�� INDr�I�"E ��NTV�E�0��+B23_Ux��=CLOWLaA�@��Q��5]FD�@@�����p�5��C($FMOS9`���В!�t23�PERCH % zCO]� �G� �C��`B2���f^c5Hi 	`��A�"UL�T ����%E��`J[VvFgTRKAqAY�� S���Q�"�U�S�q8���2QpMOM��	�@��Ȁ�����#���S�]#�b�DU���"S�_BCKLSH_C�"e���F]��3���;d�2Fj�1CLA�L�`#Bő�PpxeC�HKQ�!uS�0RT�Y��8�D�u���_�Ws�D_UM���fCณ�!��c$0LMTk�_L̀Y�dm�wE}"p{ p%u(`��%Rct XPC�AB XH�p��%�eCP��z��`�'CN_ �N�`��vm�SF��IV c2�aG��q�"��x7CAT�nSH]� � �$�6��aF��+!��̎ � PA�d�2_P�e�S_���`�V�@���S���eJG!�[����K@OG�w�RTORQUU0���C�Y� �0�B�Q� �_W�U�T���8��7��7�I*?�IM�I�F'�*������ VC�0�����1��W�ǟ���JRKל��떷�KDB� M�ӷ�M���_DL�6RGRV�>�7��7���H_p���^ e�COSr�s r�LN����ڕ�� ���� ��i�Ӫ����b�Z���F�MY����~�@ᆫ2�THE{T0fENK23��\����CBa�CB�C��AS����i�0�����a�SB���Nl�GTS��$1Cr����}���У$DU�`?W����1�������QQ��ws�QN	E��y�I���c}	M	$P�AT�}ņ�d�o�o�LPHr�[�5E[�Sڕ������Х[ ߦ������V��V��ȑ��V��V��V���V��V��V�V�H��A־Ҷ�;��ت��H��H��H��H��H�O��O��OTJ��O��O��O��UO��O��O�O���F[��������S�PBALANCEl��qLEɰH_T�SP��5���5�ЦPFULC9�`�H��`�Х"1�mUT�O_�`ȅT1T2���2N�a�-@����Qb�@�1"��QT�LPOV �(�INSsEG�AREV���@ADIFuUG1ٙ,s1�	@OB"haA��W2�-@�a~ �LCHWAR2�AB���U$MECH��!��1��fAX�QPFt�vǂ�� 
���E7ROB�@CR�"���r�DO_�DAT�� < �0�O1�by1s�{BE$ON!CD_d@y0 �0`u` �� %�0�T@A�aT#x2L̀@�`CKx2� CT1  %�`�!N�@��8�@R3`y1������ MP��3E5 $I�R���1�`�/PN2MCAI��1�2%_]C#/ !�0R,��COD7FU�0FwLAGx2ID_O`�V% ��G_SU;FFi� �0�14 �1�DO� �O�(GR]��$ ��$��%��%��$^  2�&HV �_FI-9
3O{RDA  �MMY36Jr2q!��$ZDT]% �	�c�4 =*.L_NAM�|d2�DEF_It80d2��4�ST��P���3��5�ISD��`0S���3R�~4�)34�q�]r�2D��b)D7D���O�/LOCKEn��#����1�"� UM�%d2�$�3�$ �5�$B�"�C�%�3�$ �4�"Q��5�D�1�#�  ���%d2�%�3�#�G:U�(gPT �4w�1Y��WuHtUC	��TE_Q� ��ZRULOMB_t�R�W0�BVIS��WITY�BA��O��QFRI���SU SI�1�QE�R��W�r�W3�Bn�$W�X!W�[(��V��_Ei�!'EAS._cSÁ�A��GT7� h M�TEW F7ZuCOEFF_O����d�\ GF�hcSU ���b�.x��$�`��C�- cG�RD� � � �$@��9XvTM^GtkE�sC,|B�ER  TTDS40�  ��LL�$���A3SV.D~x$�V0q��}d0� rSETU�2c2 �� � �p� "@ID�r��qCAD�vi2�CA_A@D��b'a�"��<@�
A;@"�2�W . R��0�q!bSKy_��c� P&T1_USER���N�t�o �t���VE�L�t�o �����I\=0���MTgC��>k��  �4 }O�NORESJ�ۂ�p ʂ� 4�"��r�R"�XYZx�#����DEBU��_��_ERR�! ,�PpeF �c7��Q`����`BUF�INDX�a��M�OR�d� H&CU7�L���'!<1��< 1$� ��A�1�O1��3�G�b�� � $SI�MUL+`F 	x�V�O�H�OBJE<S��ADJU�b�F��AY�0��D%��OU0���r!2=��T��T���S�DIRX�`�/ =��`DYN7b�b��	T�y�R�QwAw¿�OPWOR^� ��,�`SYSsBUm��SOPޡHZ��q�U�/ P@���PAw��q��V�OP� Uw��T+!A@�IMAGbJ�&C��2IM���f�INE`7�e�RGOVRD�� �x�B�PD�d��`S�*P/C����Li@B4���qP�MC_EE0Z�ANbm�M�!A*219 A7����SLS�k��� �� OVSL:SiRDEXA�0"&�2���a_��>� � ��>�� H�]�Xșb�}�C� f0��Z��q�¹sj�� @��4���O^ RI�� ����* �������`��PL�  _$FREEȂEıQ�a1�Lj����yT� h ATUS�p$TRC_T|�i�@�BpJ�3��tCp A�E0k�� D& @�)�=Ҧ��>�1�`J���XED��u�Ҭ��wԳð��r�C�UP�@�1PX�j�=��D3�s���Gȅ�>֠$SUB2����A2���JMPWA�IT��M�J�LOW�
���$RCV!F"!��M�Rq�ɀ�CC��R�����IGNR_PL��/DBTBh P�1�#BWB ���UY���IG'����� TNLN����R��dB�PyN� �PEED��>/�HADOWh ���E.�>�=��0�SP�� � L�&� �1^�
�l�UN!IE�n�y���R�ЗãLY:0��<�/�P4��j��>�$�D���L��NPA�R@T���*���P��k���bARSIAZG$0 3�1�O� ~�ORMATT¡p��S��MEM�(��UX͠��O1sPL[ Ʉ� $Ӂ~^QSWITCH�Z�aW�AS��P��QaPLB AL_� �y i�OPBԱ�PC�D�qP���J3D�� T�`PDCKͰ�2��CO_J3 PH��BE��a������b��˰ �� ��PAYLOYA�S_1Z2Z� J3AR��yfx�u��TIA4�u5�6�MOM @�����ŀBa��AD�����PUB��R�!%�!%����kg��` I$PI���U���_Xr*��]Zr*I
+I�+I�#�VA�& ��&������8}���"�HIG�"� b�[�6[�b��q�6�K3$8��39��b�SAMP�Њ��47�3b�'MOVU���,��1 ��@���4 ��6[�g �9u��������5RaN2�5INLR`k3H 9KDb�J_H6D_KK/GAMMESF��$GET}�f��iDC��
�aIB�b:�I'�$HI�TaALР��FE��X�P�L�PVLW�M<V3\�Y`VV�b�&��C���CHK���� ��I_j0.a���T QaE�W���&�Y�� �$� �1���I�pRCH�_D~���Ѓ�HpL�E������Uh?`���MSWFL��M.�SCR��7?��f`�!�e ���P SVt�Pxpm��g�a�w{pSAV��t�e/�NOCC��0�D�` �DS}![ᡑ)[� �[zK{� �%�xuD 3�y0�B��6�7�2�� 8�6�K8�w�u�s��10�T�L4`g�� 7� �SYLq#V�
G��SU�����>� ��*�V��SJ�V�q��`$�� �Wp����A Ȋ��� �M̐��CL �������h1 �M �M�aU"� � 9$5�Ѵ$W���� P�T������"�� )��������A�@�ųX@X��O*WAZp��M ��� ��QOM�S]0BT8fx�CONHb��tiC_s� |� ���`�H��H���`��u�`����E Q��*��b���z�,�P�PMW�Q}U�0 � 8���QCOU�Q0QT�H��HO7��HY�S/ ES�1�UE�ޠ�b��O ��  b{ P܀�E��UNE��j�V�O2u � �Py�=����a���ROOGRAX�I�2��O��<�ITK`�� ��INFO��� �{p���I���OI� (ԀSLE�Q��۱�%۰s�ױS�_EDO�u � �����K�1��QE�PNU+�%�AUT<
q(�COPY�10(I� �pM�ANS�W�^�VPRUT� Z��NFE�U�$G�A������PR�� ~�� � �� |����<�US�R_TS8���TP���KLNA�4CLl��%�TP$ֿOPTION��G t�>��"R�R�S��Rל���LD@�� ?�� |���A���z���M��PA�S���P���PRG_�(Ҟю�6��= ���e�  �PI���CH� �����8/�!��_OVbqh/����M��PT1�T�W�STATU2#I����AP� ��MO_WA����X����S�P��w��P�CR�C���aS䀜�]�p��T�f�x�������� ,��H	Ep"p�Ai�h!U k�~�� 1� ���KTܥ� < �N�TRIE#SmEݠNC�� a��j�Q�BѠe��Q�������G��LU��PRI�������WRK��� ���SV���ܢ�&Sx2����EXEC��yR鰌� �t�@1���(�:�$��`~T � Ơ�ELE�2� ���GADJ�� 5h9�X��MI=c��(����W�P�c`��3� R�EXT_�CYC*��RG�N��$��,���L�GO�S�NYQ_	Fu 8"Wj@�V����C`aLAKc���`�����@���PIF�!{�$��_GKc���2�Mk��2�q!W`�LAST!�qb���� �z�ENAyB*��EASIX! �r�2��P�G"��ay& �@�@�S�?a�����Zc�"ABCѤpE䀰"0V;!�&BASq�&�B]�U@0�@p�$�!�'RMS_TR�#WAH`3z�SP��4!�$
�d���7�	��  ECg�3Dk62j792ۀ��pn�2�7��MfDOaU2�Cd��bPR�zm��GRID��C�BARS�&��Y#$��� O���һ`.�D��'�!+BO��.i� ���L#0���R��<A�YESRV�(�)ZDRFDIpT_� t@�D�`�G� �GT�АG5�I6�I7�II8rAF��m�+�?$VALU�#�e�k$�p��Fh�� ��U$q}�$C*��h|�AN�cR !�ъQ�qTOTA�#� �vRPW}I�1�TR�EGEN�Z�R��X�8Q�t庡@V٠TR�#"�Q_S�`�W�P��#V��b��!E� #�0���r<�?�RSV_H�0DAٓ`P`GS_Yqz��S�{ARِ2� �IK�E��PRB0%_�@�+dhD�A�5� �4��?�&�[�hSL9G�`�� @\�P� ���݂p� Sy�1$DEqAUO�2�װ�`�TEr�m�� �!�Q���J�fQ�C��IL_M�~pV�"|Л�TQ٠�ӓ�R0C��m�V�{C�}�P_}p� �sM�yV�1�zV1�{2�{2��{3�{3�{4�{4 �zo�� o2o�w�s��vp2IN��VIB�T�t��2��2��2��U3��3��4��4�����rIqf����D $MC_F��|	���xfSM����7�+��3 �9��5q� KE�EP_HNADD"$�!f�� p�C��(�A��A%�����Oҡ e���#�`������RE|�r��!��Õ�ڑߘU$�e��HP�WD  f�S�B��+@COLLAABt9PpgQ������O�r��N3ڞ\�$FLj0�!O$SYN�t�M;0�C�b��PUP_D�LY��+�DEL�A��!{�Y�pAD�RaM�QSKIP�e�� ���>�OR`f�|��1Р�RRg� �o�j2����w� �������@��@���@��@�9�!��J2RG���bEeX� T���ITS���;�b����ab��`RsDCKQh�� ��R-1TOR��pp1�R����!0 �m4R�GEA�R û2F�LG� �W�L�m4S�PCĲ�嵰ds2TH2N0�������  ��0POwS11W�� lW�`��)r��U#J�AT���CH�UjTns��I�N����m4��TO<�o2HOME��ʠ
��2���ϸ�����P�� �^��3���#�@5�G�Y�k�}��4���߲��������ߏ�5����/�A�S�e�w� ��6��䀚����������7���)�;�M�_�q�W ��8���@�����������S*�
���,1�óPJ��=!ڒEh��`0Y��lV�IOaq�	�IO C0̡R�WE��� � s�ӱq���PgS �n�$DSB��;"�eS��C��C0�S2;32�� ���y��5pICEU�"澠PE��i!PARsITRadQOPBR��h"FLOW�`TR`k qR��0i!CU�=Mh#UXTA+�i!�INTERFACpl"_��SCHSq� tW� �00�aT�3$� 1`OMj`s�A/�<0I$�� �0ADn�� T� aCS X��85(#[pEFA�p^��[�RSP�Sq���Zp$USA�w��q"	�EX�I�O��: �PY�%&_`�r9Q� �&WR,��7I
�0�(�MFR�IENDM1<�$�UFRAM�d0TwOOL$6MYH ��2LENGTH_VTE
4I�qM3�0�$SE:[9UFWINVQ@S����RG�2�0ITI��T7X|�e7�6G2�'G1A��#�2�72�`_2o�O_jK  <�=1�p'�>�Ce#ju�Cn�b2�1&F �G&��Sq�r�j�5�J�(�c�b�����g$�X � E_MY CT�#Hа�(���$e#%Gn�W� �G�B�D=DĠLOCK�E��`�a�AT0�$?F 2�W��!��)�1�(�2�+2O[3�+3�*?Y�Q�)]Y�Q�M� c� cVp�@��U@�9FBTp����(S*���F�"k @2��A�5�E��Nb�a3�}1`4ACdiP!Rϰgf}E�SS@����P�m c$M� 0�0�F4Pﲰ�T4PA�W�e �0��
b%�S��� �	aR�3!`r�q$RUNMN� AX�@A0�LH1��rTHIC��!�Ӡ4%�FEgREN�auIF���#qI�'gsM�`G�1�h�tL �y�o n�v_JF�wPR@����RV_DATA�� ��̐��- ��AL� o�v�� ���q  ?2� �S�O?�	� �$Ű��=s�GROUǱ7��TOTt7�DSP>N�JOGLI�y0'E_P���O.q��� @�K. _MI�Rj����0M�B��A	P�AiAE� ˀ5$t��SYS���t�PG���BRKB4&��A;XI]  ��#��9�`A:�C���B�SOCB�� N>�D�UMMY160��$SVU�DE_O�P�SFSPD_�OVR�`�p1�DLy�|�OR��/ N% b��FNq��g�OVj�CSF��p���BFٖ�����3�.1�LC�H����RECOV(x�� g�W��Mg�/�Fj�RO�J�v�_p�p @Y0VE�R�`� OFS�0C�p3WD��+���J�X�"ąd�TR���аE_FDOĆMOB_CMǱ��BZ��BLb��Ѣa�dV@BA�R  O`���Gҧ�AM�Š `�R�-�_M頷P��_�OT$CA]�P�D�d�HBK$!3&y��IO�%����APPA|���������8���_�DVC_DB �3�4!�;��ő1	�R��3	�X�ATIO��x�qU�#\��CABs� �"�3�@<�i@��Qg��_�3&SUBCP	Ut�SR@	�����% �S���S��~�$HW_C�S���%SA�1�p�$U�NIT���A�TTRIӀ"�t�C�YCL�NECA�Nµ�FLTR_2_FIt3T�%�Q�LP��_p^p_SCmTCF_�F_܌��*�FS$��CHA�!�������RSD\� +�>sv� _T�PRO:�,���EMe _G��9T���Q ���Q�U�DI� 5$RAI�LAC��YBM �L!O.�@3V��aJaX�XSaX�R�PR�S(AI�`��Cݱ_	Q��FUNC}�`bRI�NG@Q!j���RA��B d�	� �r�	�WAR�se�BL"A�:�A3�/�6�/�DA�
�t�:�3�LD l��A��q�Ja��TIRb��2�v�p$h RIA�V.AF��P�����J���\PR��p�MO9IЬ�DF_F0�l!!�LM��FAY0�HRDY�$ORG���H�A!|�;MULSEF0Ӄ���QV�J��J�������FAN_ALML�V��WRN�HARD� $&�@@@�B�2��/��_&��3&AU�R�ԸTO_SBR߲$[��/�߳��GMPINFp$�Z��e7REG�&NV" �#f�DA10��FL��}�$Ml�_u�R�2�p�����t��"�� �0
1$.�!$Z'q���#��� �؃EaGR`7�l�'!ARI��]�T�2��6%`��A�XEQ�ROBN�RKEDN�W�1�_�-�0�SY	�a!��&S��'WRIY0:&��SCTRM�%���Eё�pC$�a@B�� ^��&5��>�OT�Ou�pJ�ARY�N�02��>��q�FI��$LINK(*$qP1�Q_�#^��B%6^�x1XYZt��:7�6OFFf�RO2w2k840BL�����4;�5����3F�I=��7�ao�d���f�_Jy��r��\3�A�� 4;8^��ATB�&Ay^BCd�ԆDUt|�A&9��TUR� !X��E>1UX� l�FGFL�P�m�4 �@ę5�)3�`� t� +1��pKs�M��T��3�Q���Rb�ǎ�ORQ2�[���H]�K` 뀚p, SaeUӃY��NzTOVE�Q'rM�� �q��U#�U"�V�  �X��WИT�u���� ��(q�Q���P
q�U��Q�W$e#$e�S[�E)Rx��	��E� ��$��bdAa�p�5�`-�<7{�x�{�AX;� �r{�)���Q2�e]��i ��i0�j 0�j�0�j@�0�jW@�j�@�j1�@ �fg �ig �ig �ig  �ig yg yg $yg �4yg DyaqUyDEBU��$���U��{�s2AB{�y���{S9Vn��� 
 �� <aH���T���T�1T�  1T��1T��1T�WAT���A��c@���R�3LA�B�2FU���GR�Og�FB�W�B_ ;�If�$���0,��1�pGU-�9�ANDP���WdX�|5Zav�  W�a{1��l�Z�{0�NT� /���VEL`A��TƑy�Ζ�$���ASS  ������mPmP ��k�SIL �]�����Ie�x|���AAVM� �K 2 0�� 0  G�5��g�s�d�.�� ��	����ͯmP1������ߦ�����(���.�c�u��}�A�BStQ  1��� <Q�¿Կ���
�� .�@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖߨߺ��� ������&�8�J�\� n����������� ���"�4�F�X�j�|� ������������ݐ$ �g �����  d��IN����PRE_EXE!C &T��0�A��IOCNVEB �Pk]@����wIO_p  1N�P $>����2��1�?������  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o �o�o�o�o�o0 BTfx���� �����,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z��������¿Խ��LARMRECOV Z���&�LMDG K�� ��,�?_IF � ���ϓϥϷ���o��������/�, 
 /�X����~ߐ���ߴ���ANGTO�L  Z
 	 A   ������PPINFO 6� 5�8�J�\�n���  B�p�� ����������!�@�E�/�U�{�h��� ����������%�7I[m��PP�LICATION� ?����h�LR �Handling�Tool � �
V9.10P/�03��
88g340��
F0�951����7DF1� ���None�F{RA� 6%��_ACTIVE��  ���  ~�UTOMOD��:��ӪCHGAoPONL� ��OUPLED 1^�� * ./@/�R/�CUREQ �1	^�  T\)
\,\,	�/�%� �$��\"���$H�%-"�*HTTHKY�/
��$\�/�/X?"? �/F?d?j?|?�?�?�? �?�?�?�?TOO0OBO `OfOxO�O�O�O�O�O �O�OP__,_>_\_b_ t_�_�_�_�_�_�_�_ Loo(o:oXo^opo�o �o�o�o�o�o�oH $6TZl~�� ����D�� �2� P�V�h�z������� ԏ�@�
��.�L�R� d�v���������П� <���*�H�N�`�r� ��������̯ޯ8�� �&�D�J�\�n����� ����ȿڿ4����"� @�F�X�j�|ώϠ��#�n%TO�й�DO_CLEAN�|�1�NM  �� \/ߑߣߵ����b.DSPDRY�R8ߪHI�[�@ l�3�E�W�i�{�������������MAX� ����!	')��X�(%"(�PL�UGG �%#�P�RC��BY�]��"����O�����SEGF�K������ Y�k�3EWi{����LAP�#�#� ��);M_�q����TOT�ALK�t�#USE+NU + ��/��"n RGDISPWMMC��;1C��&;�@@�$O�0����#_STRI�NG 1
�
��M�S��
~!_ITEM1�&  n��/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�?��?I/O S�IGNAL�%�Tryout M�ode�%Inp�:@Simulat{ed�!OutLLOVERR� = 100�"In cycl@E��!Prog A�borVC�!6DS�tatus�#	H�eartbeat��'MH Fauyl�G�CAler�I O�O__1_C_U_g_8y_�_�_ ӄ+ і/�_�_ oo$o6o HoZolo~o�o�o�o�o��o�o�o 2�_WOR���+jq�_D� �������"� 4�F�X�j�|�������8ď֏�PO�+�A ��{��1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u���	�DEV���%���ٯ ����!�3�E�W�i� {�������ÿտ������/�PALT �]V��0�~ϐϢϴ� ��������� �2�D� V�h�zߌߞ߰���D�GRI.��+��n��� "�4�F�X�j�|��� ������������0� B�T�f����R�]�� �x���������  2DVhz��������
��PREGZ�C��j| �������/ /0/B/T/f/x/�/�/��/M�$ARG_�jpD ?	�����!� � 	$F	+[8]7�G&9�� SBN_CONGFIG@�+DACB�>1CII_SA_VE  Dc1�Z2� TCELLSETUP �*�%  OME_I�OML%MOV�_H�0�?�?REP���O�&UTOBA�CK�1�)`1�FRA:\0c O0}0'`�@�0[F � �lK_0 1�8/02/09 �11:06:040'80�O�O_�OLL��'_N_`_r_�_�_�_0�<_�_�_�_ oo0o�_Tofoxo�o �o�o�oKo�o�o ,>�obt���������  GA_�*C_\ATBCK?CTL.TM�����1�C�U�KINI�Y�0V5$CMESSAGr0|�}1|� ��ODE_D�0u6V5f1��O����$CoPAUS�!��+� ,,		� '0�%�,��L�6�X� Z�l�����ʟ��Ɵ �`�$�� �Z����~��TSK  �x[Oa�'@UPDT���z�dˠˆXWZD_ENBz�R:Ԧ�STAy��!˥�!X�ISD0UNT 2��%c1|0� 	� N{� ��%���T���� ��(06��D��W�^5�V���0^��  �v  6e����o��ڿ��׿���MET��2��~3� P5�@��rA�1͹A��6�33A8�@��ߠS�6��^�8�8R32�4�5�7�A��6���SCRDCFG 1�%;=A �z5z2��������	��-�TO0Qv9��}ߏߡ� ������>���b��1� C�U�g�y�����'*A�GR���ߏ���pN5A�0�+	*D��_EDx�1��� 
 �%-�pEDT-���:6�Z�����~E �+B)�0�'2_�6"���  ����2���;��& �t���_����N����3��+=�@+r����4c ���=��>P�t��5//�|/� =X/�/
//�/@/��6�/k/H?�/=$?�? �/�/~??��7�?7? O[?=�?[O�?�?JO��?��8�O;��O_�� >�O'_nO�O_�O��!9__�O�_�O�>�_��_:_L_�_p_��CR ��Owo�o8MRo�oo�o�o:o���NO_�DEL����GE_�UNUSE����I�GALLOW 1���   (�*SYSTEM�*�	$SER�V_GR�{wp��REG�u$�s�wp�NUM�z�s�}P�MU#p�LA�Y/��PM�PALy��uCYC10~���=�ULSU��}����sLS���BOX�ORI�uCUR_�y��}PMCNV6�vy�10-�߀T4DLI`�w��t�	*PROGRA�tPG_MI�/�A�AL`�T��p�A�Bl�w~$FLUI_RESU�(���L��l�o� ��(�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�l�~����� ��ƿؿ���� �2���h��LAL_OU�T f{����W?D_ABOR�G~����ITR_RT/N  �T�Py��?NONSTO����� ��CCG_C�ONFIG  ��L������&�8���E_RIA_IDp���`�Tq��F?CFG ����]i�_PA��G�P 1s�����������߾�C��P �"���C��Ce "�("�-�C8"�e@"�H"���CX"�U`"�h"�p"�x�U�"�"�"�"���������U?����HE�`ӥ���G�_P��1��  5�s6�$�6�H�Z�l��~���B�HKPAU�S��1��`�  -����������� B(fx^��������,>�O�m�s��WXpCO�LLECT_m�Ƨ���uEN����Or�NNDE�}����b�1234567890��R�q����F�S
 U�]��Q)0/ U/�l//A/�/�ks/�/ �/�/�/�/&?�/?? n?9?K?]?�?�?�?�? �?�?�?�?FOO#O5O �OYOkO}O�O�O��q;2� ��IO  ���X���X_j_|_�_&WTR���2!
]E� AY
�O�^�"5]�ZHu^�_MORR#��� ���Oe 	  OigoUo�oyo�o�k(bT��Q$6m,Hu?����sKPKtKQARJ��PR&�g��Xj|�
I�k ����Q��rZӝ�u� �a�PDB�T(���Dcpmidbg�T��f�:��N;�p@���d�_  ��N>�ݏ��ܺ���%�����mg�o�:����f^������@ud1:ܟ��Z�?DEF '@S�)�c�buf.txt�^����_MC/c)��Sd����.d*��u���ѥ>�vCz  B*!�`�Bΰ�Cy�CCI;�p����C򠧺z�`DD�4VD��D��J0?M�D��I�DD.a
�F��F��F�U�CH�J�F2�y�b�a��
�g,
\T�k!KPU�`KP�`��`ɐ�T�m�`E��@ D1�D�  �E	� D�@ �˱2�| Fp� F"� G=��fF��G'i�
�G>�Gg�� GK  H��<=H�&H�yMZ��  >�?33  `C���1n���r�5YKşb�Q�Aq�t=L��<#�eMQ���Ş�|�RSMOFST� %/�:HP_�T1��DE -�*���Qw�KQ;壍��ϩ�?��Ϛ<�2��ES�T)�+/���R.XX��զC4y��z	�KPm�{����T��B�R��p����?�KP:d�
��T�_)�PROG ��Ʃ�%o�I��.PN�USER����\�K�EY_TBL  �����h9��	
��� !"#$�%&'()*+,�-./�:;<=�>?@ABC)�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������#��͓���������������������������������耇�����������������������A�LC�Kg��^�g�STA�T����_AUTO�_DO�����I#ND���tR������T2*z�STO��NTRL�L�ETE�q
_S�CREEN ~6jkcsc��Ub MMENU {1/%� <8� 7���u�=̓ @yPb���� ���-///c/:/ L/�/p/�/�/�/�/�/ ?�/ ?M?$?6?\?�? l?~?�?�?�?O�?�? OIO O2OOVOhO�O �O�O�O�O�O�O3_
_ _i_@_R_x_�_�_�_ �_�_�_o�_o,oeo <oNo�oro�o�o�o�o �o�oO&8� \n�����ƙ��_MANUAL�f�DBCO R�IG���&�_ER�RL%�0��X��Eߖ����� C�NOUMLI2�M������DBPXWO_RK 11������,�>�P�b�v�DBwTB_| 2r��ѣ��ؤ	�DB__AWAYK�X�/GCP ��=<ж��_AL2�����G�Y�e ���<�_e� 1}3� , 
	�`G���5�r�|�_M �I��Ĝ@|���ON�TIM����ɼ���
v��MO�TNEN��m��R�ECORD 19Α� �z���G�O�B�0���Œn��� ����;���ӿB���f� �-�?�ֿ�u�俙� Ͻ������ώ�߆� ;ߪ�_�q߃ߕ�߹� (���L���%�7�� [�����ߣ������ H���l����E�W�i� {�������2����� ��A,:w�� ���.��d �=Oa�p� �*��/��9/ �]/��/�/�/�/R/ �/J/�/n/#?5?G?Y?��/��TOLERE�NCÔB��ѐL���C�CSS_C�NSTCY 2:J�����\?
���? �?�?�?OO,O>OTO bOtO�O�O�O�O�O�O��O__�4DEVI�CE 2;�; ��i_h_�_�_�_�_��_�_�_oo{��3HNDGD <�;�7�Cz7nLS 2=P]/o�o�o�o�o��o�o1o�2PARAM >#��u\��4SLAVE �?Pm<g_CFG� @9sd�MC:\�0L%0?4d.CSV
��c�	��"A �sC	H�pbab�~�-�
vW�v�J�Z�H�<G���JP�z�o_�
�����~tRC_?OUT AP]���_SGN B���&j���27-FEB-18 10:35�p��09�1:�06�pyV LIX�9�5�~6����+��i�Þ�����I�|uVE�RSION ���V4.1.�0��EFLOGI�C 1C�; 	r��ԙ�䝶��PROG_ENB���Xf�ULS�� �Wf��_ACCL{IM���ss��C�WRSTJN`��٥����MO����ur��INIT cD�:�� ��wOPT`p ?	�����
 	R5�75s�74�6J��7��5���1��2��r�B���ѤTO�  ݭL�����V.��DEXp�d{������PATH {�A\������s;HCP_CLN�TID ?��qs� ��3N�}1I�AG_GRP 2�I�y ��� 	 @K��@G�?����?l��>����dʘ��1��d������0����?�b�?�� �i�^?�V�m?Sݘd��f403 6789012345>�ܓ���� ��s���@nȴ@i��#@d�/@_��w@Z~�@U/�@O�@I��@D(�d�\О��@��tp�p�ѓ0Ae�0�0�pB4d̡]Pd�ݨ��
[�1���-@)hs�@$��@ bN�@��@e����@�D@+���ߦ߸Խ��������R��@N�@I�@D��@>�y@9���@4��.v�@(��@"�\��%�7�I�[���L��@Gl�@BJ�@<z�@6e�0��`@*y�$�?�@�������������=q@�q��F@|��@33@��R@-?����?��`?�++�=�O�a�s������-@&��@�}��!�?�?� � �����������׋� ������C !Sy_�� ��	/�/Ţ��p�@�ш���, ����t!Y����?��z�!��5AF��!4�� ��L4�R�!��@�p]��"�Q��"-� �� Q�@�U ��Ah���=H�9=Ƨ�=�^5=�0��>���o=�,'?�,7�� ���C��<(;�UC� 4�¤��k?��d�A@��? ��3/�?;-�?�?�?�� d4�?)O�?9O_OAO�O��O?)>��y�B��R=���=���z�A�ͽ�G��OG����u�uWW��.T@�pғ6�̷�uB���X B��B��B%C��͟��_p^'Q�©U���Q�Q�L䏁\c����*���� B��@B��B��A��@���_c�0o��< ~�5o^opo?�o�oo��ot[�o�bd�D����:B����C�з��B���?� �o3�oWB{f��d�v�CT_CON�FIG J��|��/�eg���u�STBF_TTSp�
��s��O�F�:���MAUj��~�MSW_CF�p�K��  ��ڊOCoVIEW"�Lb�����Lo��Ə؏� ���S���7�I�[�m� ��� ���ǟٟ��� ���3�E�W�i�{��� ��.�ïկ����� ��A�S�e�w�����*� ��ѿ�����+Ϻ� O�a�sυϗϩ�8����������'�s�RC[�M�/�!��5�_� �߃߸ߧ����� ���SBL_FAUL�T NR�w��G�PMSK�-��pTDIAG O�yچQ'��'��UD1: 6789012345���r~��w5�P����� ����� �2�D�V�h� z���������������z�5ِ2
��.�vTORECPc�u�
�� u��6����� �/ASew �������
�/x�UMP_OP�TION�&�3!T�R[��*�T%PM�E�G/Y_TEM�P  È�3�B�P� ��Q�$U�NI@���!O�YN_BRK P��~R�EDITOR9!�?!�/�"_K ENT� 1QR�  �,&PROG_�1 -!/{m&-?BCKEDT<?N?�ߝ?�r��?�?�? �?�?�?"O	OFO-OjO |OcO�O�O�O�O�O�O �O___T_;_x___ �_�_�_�_�_�_o�_ ,ooPoboIo�omg� �MGDI_STA��%�q�!�%NC�c1Rb� ���o�o
".
".d	/L^p ������� � �$�6�H�Z�l�~��� ����Əa%ݏ��� !�9q!�G�Y�k�}��� ����şן����� 1�C�U�g�y������� )�֏����0�:� L�^�p���������ʿ ܿ� ��$�6�H�Z� l�~ϐϢϴ�ί���� ���(�2�D�V�h�z� �ߞ߰���������
� �.�@�R�d�v��� ���ϴ������ �� <�N�`�r��������� ������&8J \n�������� ���*�4FXj |������� //0/B/T/f/x/�/ �/���/�/�/?" ,?>?P?b?t?�?�?�? �?�?�?�?OO(O:O LO^OpO�O�O�O�/�O �O�O _?$_6_H_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�O�o�o�o�o_ .@Rdv�� �������*� <�N�`�r������o�� ̏ޏ��
&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφ� ��� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~��ϴ������� �� �2�D�V�h�z� ��������������
 .@Rdv��� �������* <N`r���� ���//&/8/J/ \/n/�/���/�/�/ �/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�/ �/�O�O�O�O�/__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�O�o�o�o �o�O $6HZ l~������ �� �2�D�V�h�z� �o����ԏ�o��
� �.�@�R�d�v����� ����П�����*� <�N�`�r���~����� ̯�����&�8�J� \�n���������ȿڿ ����"�4�F�X�j� �����ϲ�������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b��ώϘ�� ����������(�:� L�^�p����������� ���� $6HZ l�������� � 2DVhz �������
/ /./@/R/d/~l/�/ �/�/��/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \Ov/�/�O�O�OlO�/ �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTonO�O�o �o�o�o�O�o�o ,>Pbt��� ������(�:� L�^�xo���������o ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�p�z� ������ʏ�����
� �.�@�R�d�v����� ����п�����*� <�N�h�ZτϖϨ�¯ ԯ������&�8�J� \�n߀ߒߤ߶����� �����"�4�F�`�r� |������������ ��0�B�T�f�x��� ������������ ,>��j�t��� �����(: L^p����� �� //$/6/H/b l/~/�/�/��/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OZ/HOvO�O�O �/�O�O�O�O__*_ <_N_`_r_�_�_�_�_ �_�_�_oo&o8oRO� �$ENETM�ODE 1S�E��  
b@b@]Eo�ka`�RROR_PRO/G %nj%\F�o��i�eTABLE  nk�O 2D�Rw�bSEV_NU�M }b  ��xatp�a_AU�TO_ENB  q�evc�d_NO�q� Tnk�asr�  *��p��p��p��pp+�p��<	��tFLTR��v�HISps`Av`�{_�ALM 1Unk� �]D�|\@+ 
�����ɏۏ�����_ir�p  nk��q�bD�a`TCP_�VER !nj!��o�$EXTLO�G_REQE�蜜y��SIZ����SkTK���u����TOL  `AD�zM��A ��_BWD$���)�%��bv�DI� V�E�)��d`A*�S�TEP;�M�a`g�O�P_DOޟ_aFD�R_GRP 1Wni/�d 	?�ܯ�`�͠n&����c?��$,�MT� ��$ ����ͣ"� 3��V�A�z�e������¿���������A�W�As�Y>�(��#�b@
 E��`B@�Kϗh>����ϲϝ�����A@�:���@�33@���Ӽ�@��߻�xD�V�͠F@ l��`�`�l�\ބL�F�Z!D�`�D��� BT��@����4�?�  ���Z�6��������5�Zf5��ES��4ݺ@��ƿ�� .b��a�XV,�����k�FEATURE �X�E%��a�LR Hand�lingTool� ^�`BEng�lish Dictionarya��4D StS�ar�d^�`�Analo�g I/O���g�le Shift���uto Sof�tware Up�date��mat�ic Backu�p_��groun?d EditW�a�Camera��F���Common �calib UI�8�D�n�O�Monoitor\�tr\�?Reliab��`��DHCP9�^�Da�ta Acqui�sk��iagno�s����ocum�ent View�ew��ual C�heck Saf�etyW�d�hanGcedW�`�-s  �Fr0�b�xt. oDIO g�fi���\end1 Err�v�L��xPsw	r��g  �^�FCT�N Menu v|���TP In� �fac�c�G�p� Mask Ex�c- gYHT� Proxy Sv�igh-Spe1 Ski���k �mmunic��onsVur� � ������connecwt 2�ncr� �struu�_�KA�REL Cmd.� Lua�R�un-TiX Enyv�� el + ��s��S/Wa�License � �Book(Sys�tem)^�MAC�ROs,M/Of'fse��T%Hk �����Y MRp�l���M�����l Mec_hStop+t�D��T%i����&x1 ئ����.od��wiGtch?�#��.y&4;OptmF?�#,�fi�.�&g�T%ulti-T"�_�PCM fun�:�9a� tiz�8�7�o��RegiI r,q�6ri��F�;F���Num Sel��%/IV  Adju�a*NWA��hMtat�uA�O��c�RDM� Robotr�s�cove{�Eem�� kn��E�BSe�rvok !0`�SN�PX b"��SN�� Cli��#^��LGibrz�C_S� �$�UPVo. t� ss#ag�5d�X� ��l!̕�X�/I��UMI�LIB�_�RP F�irm��^P�A�cc�!�TPTX���Telnl �_�Qx[�h%�]orqu��imulau�6�U���B3&+ev.̜U��ri 8oUnexcept1 ��@n�eQ��VC"S�rlc�(V��r� o*uU[${S6PSC�2e\SUI��Web Pl�F�~Q��t3+��ZDT� Applj^�i�P� a<Y� Gr{id�Aplay�(�P��Rr.��X����1"� ��200yi���scii+�VBLoad  ��U�pl;���Pat)6(�yc���@�` �RL�V �y~ MI Dev$ � (QM"�6��7s�swo���/64MB DRAM�Β�FRO��-�ell��B�sh̑؟�1ce;���pa
!��sty��sAB��t�^0.���@k����6� 2�a��poCrt?�@ R��q$�T1p�	[� ��d�N'o m�@{�c�d�;OL[�Sup��}1HOPT �,�Z�9S� cro�L�C�UUL��NF���ues�tUS[�e�te�xqdUp��_PqP� %OTou(0P+�s{rt�C��stdpn�ks� �SWIMEST Mfv�F0]�b��W� �i�{Ϩϟϱ����� �����7�A�n�e� wߤߛ߭�������� ��3�=�j�a�s�� ������������ /�9�f�]�o������� ��������+5 bYk����� ��'1^U g������ / �	/#/-/Z/Q/c/�/ �/�/�/�/�/�/�/? ?)?V?M?_?�?�?�? �?�?�?�?�?OO%O ROIO[O�OO�O�O�O �O�O�O�O_!_N_E_ W_�_{_�_�_�_�_�_ �_�_ooJoAoSo�o wo�o�o�o�o�o�o�o F=O|s� �������� B�9�K�x�o������� ���ۏ���>�5� G�t�k�}��������� ן���:�1�C�p� g�y�������ܯӯ� ��	�6�-�?�l�c�u� ������ؿϿ���� 2�)�;�h�_�qϞϕ� �����������.�%� 7�d�[�mߚߑߣ��� ��������*�!�3�`� W�i���������� ����&��/�\�S�e� ���������������� "+XOa�� ������ 'TK]���� ����//#/P/ G/Y/�/}/�/�/�/�/ �/�/???L?C?U? �?y?�?�?�?�?�?�? O	OOHO?OQO~OuO �O�O�O�O�O�O__ _D_;_M_z_q_�_�_ �_�_�_�_
ooo@o 7oIovomoo�o�o�o �o�o�o<3E ri{����� ���8�/�A�n�e� w�������Ǐя���� �4�+�=�j�a�s��� ����ß͟����0� '�9�f�]�o������� ��ɯ�����,�#�5� b�Y�k���������ſ ����(��1�^�U� gϔϋϝϷ������� ��$��-�Z�Q�cߐ� �ߙ߽߳������� � �)�V�M�_���� �����������%� R�I�[���������� ������!NE W�{����� �JAS� w������/ //F/=/O/|/s/�/ �/�/�/�/�/??? B?9?K?x?o?�?�?�? �?�?�?O�?O>O5O GOtOkO}O�O�O�O�O �O_�O_:_1_C_p_ g_y_�_�_�_�_�_ o��_	o6o-a  ?H551+cQa�2VfR782Wg5�0WeJ614WeAwTUP{f545{h�6WeVCAMWeC�UIF{g28�fN�REcf52�fR6�3bgSCHWeDO�CV�fCSUcf8�69{g0�fEIOuC�g4nfR69�f�ESET�g�gJ7ީgMASKWePR�XY�h7WfOCO�_x3�hnfgpzhyh5u3"vH�xLCH�v�OPLG�g0�vM�HCR�vS�MA]T�fMCS�h0jw{55�fMDSW[�v�wOP�wMPR�vp�`�v+pzfPCM�g�5��gp�f���51֞g51҈0�fPR�S^w69�vFRD޶fRMCNWf93�zfSNBA�g�wSHLB3�MU��`N��2zfHTC�fTMsILch"vTPA:voTPTX��EL&�t�"w8mgJ95�fwTUT�vUEC�vwUFR�fVCC
��O�VIP��CS�C��pIWeWEBn�fHTT�fR6�h�ؘCG]�IGE�I�PGS��RC��D�G�wH75�fR7�QwRЈR66�x2v�vR6UgR55�q4Vf�`VfD06�f�F(�CLI���gC�MS:vW��fSTY.�TO^�7!w�`�fwORS�R68zf�M �NOM:vOL�A�OPI��SEN�DcfL�S��ET�S��+p��CP�g7�8VfFVR:vIP=N��GeneWd2h ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߡ߳��������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻߀��������'�9��  H55�1;�U�2Z�R78�2[�50[�J61�4[�ATUP��5�45��6[�VCA�M[�CUIF��2�8��NREk�52���R63j�SCH�[�DOCV;�CS]Uk�869��0��EIOC�4z�R{69��ESET�����J7��MASK^[�PRXY��7[�OCO��3��z�����53j�HHL{CH��OPLG��0*
MHCR��S�MAT
�MCSڪ�0��55��MD�SWOPM�PR
'�

w���PCM��5i��� �Z51��51�0n��PRS��69

�FRD��RMCN�[�93��SNBA��ISHLB+*M�Y+'��2��HTC���TMILk�j�T{PA��TPTX�*�EL*� j�8y�J�95��TUT
U�EC��UFR��V�CCJ<O�
VIPN�*CSC�*X�I[�wWEB��HTT��R6�<CG�;I�G�;IPGS�:R�C�*DGH75ֺ�R7��R�R6�6*2*
R6Y�R�55zL4Z��Z�D�06��F�LCLIJ��CMS��P��STYz;TO�;7�i����ORS�
R�68��M�NOMv��OL�OPI
J�SENDk�LY;S�h\ETS
Jw�+C�P
�78Z�FVR��IPN�*Gene[�:�aoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /ASew� �������� +�=�O�a�s������� ��͏ߏ���'�9� K�]�o���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹߀��������%�7��C�STD>�LANG_�Z�r� ������������ �&�8�J�\�n����� ������������" 4FXj|��� ����0B Tfx����� ��//,/>/P/b/pt/�/�/�*RBT^�OPTN�/�/�/�/>?DPN]�-? ??Q?c?u?�?�?�?�?��?�?�?OO)O;Oted _�6�eO wO�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�o�o#5 GYk}���� �����1�C�U� g�y���������ӏ� ��	��-�?�Q�c�u� ��������ϟ��� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_�W_i_{_�_�_�_  ��_�_�_�_o o2m�999e�$FE�AT_ADD ?_	���fan`?  	6hwo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� Y�k�}�������şן �����1�C�U�g� y���������ӯ��� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_�qσϕϧ� ����������%�7� I�[�m�ߑߣߵ��� �������!�3�E�W� i�{���������� ����/�A�S�e�w� �������������� +=Oas�� �����' 9K]o���� ����/#/5/G/�Y/YdDEMO �Xfi    6h�-�/�/�/�/�/? ??A?8?J?d?n?�? �?�?�?�?�?O�?O =O4OFO`OjO�O�O�O �O�O�O_�O_9_0_ B_\_f_�_�_�_�_�_ �_�_�_o5o,o>oXo bo�o�o�o�o�o�o�o �o1(:T^� ������� � -�$�6�P�Z���~��� ����Ə����)� � 2�L�V���z������� ����%��.�H� R��v���������� ���!��*�D�N�{� r����������޿� ��&�@�J�w�nπ� �Ϥ϶��������� "�<�F�s�j�|ߩߠ� �����������8� B�o�f�x������ �������4�>�k� b�t������������� 0:g^p ������	  ,6cZl�� ����/�/(/ 2/_/V/h/�/�/�/�/ �/�/?�/
?$?.?[? R?d?�?�?�?�?�?�? �?�?O O*OWONO`O �O�O�O�O�O�O�O�O __&_S_J_\_�_�_ �_�_�_�_�_�_�_o "oOoFoXo�o|o�o�o �o�o�o�o�oK BT�x���� �����G�>�P� }�t������������ ���C�:�L�y�p� ���������ܟ�� �?�6�H�u�l�~��� �����د���;� 2�D�q�h�z������� ݿԿ� �
�7�.�@� m�d�vϣϚϬ����� �����3�*�<�i�`� rߟߖߨ��������� �/�&�8�e�\�n�� �������������+� "�4�a�X�j������� ����������'0 ]Tf����� ���#,YP b������� �//(/U/L/^/�/ �/�/�/�/�/�/�/? ?$?Q?H?Z?�?~?�? �?�?�?�?�?OO O MODOVO�OzO�O�O�O �O�O�O_
__I_@_ R__v_�_�_�_�_�_ �_oooEo<oNo{o ro�o�o�o�o�o�o A8Jwn� �������� =�4�F�s�j�|����� ��̏֏����9�0� B�o�f�x�������ȟ ҟ�����5�,�>�k� b�t�������įί�� ��1�(�:�g�^�p� ��������ʿ��� � -�$�6�c�Z�lϙϐ� �ϼ���������)� � 2�_�V�hߕߌߞ߸� ��������%��.�[� R�d�������� ����!��*�W�N�`� ���������������� &SJ\�� ������ "OFX�|�� ����///K/ B/T/�/x/�/�/�/�/ �/�/???G?>?P? }?t?�?�?�?�?�?�? OOOCO:OLOyOpO �O�O�O�O�O�O	_ _ _?_6_H_u_l_~_�_ �_�_�_�_o�_o;o 2oDoqohozo�o�o�o �o�o�o
7.@ mdv����� ���3�*�<�i�`� r�����Ï��̏���� �/�&�8�e�\�n��� ������ȟ�����+��"�4�a�X���  {�������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o0B Tfx����� ����,�>�P�b� t���������Ώ��� ��(�:�L�^�p��� ������ʟܟ� �� $�6�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�j�|������� ��������0B Tfx����� ��,>Pb t������� //(/:/L/^/p/�)  �(�!�/ �/�/�/�/�/
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O�O�O�O�O�O �O__&_8_J_\_n_ �_�_�_�_�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�o 0BTfx��� ������,�>� P�b�t���������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l�~� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� ��������*�<�N� `�r߄ߖߨߺ����� ����&�8�J�\�n� ������������� �"�4�F�X�j�|��� ������������ 0BTfx��� ����,> Pbt����� ��//(/:/L/^/ p/�/�/�/�/�/�/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�?O  O2ODOVOhOzO�O�O �O�O�O�O�O
__._ @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�o�o�o �o&8J\n �������� �"�4�F�X�j�|��� ����ď֏����� 0�B�T�f�x������� ��ҟ�����,�>� P�b�t���������ί ����(�:�L�^� p���������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ����������  �2�D�V�h�zߌߞ� ����������
��.� @�R�d�v����� ��������*�<�N� `�r������������� ��&8J\n �������� "4FXj|� ������//@0/B/T/f/x/�!� (�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| �������� �0�B�T�f�x����� ����ҏ�����,� >�P�b�t��������� Ο�����(�:�L� ^�p���������ʯܯ � ��$�6�H�Z�l� ~�������ƿؿ��� � �2�D�V�h�zό� �ϰ���������
�� .�@�R�d�v߈ߚ߬� ����������*�<� N�`�r������� ������&�8�J�\� n��������������� ��"4FXj| ������� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟������0�B�T�f�x�����$FEAT_DEMOIN  �����������I�NDEX��������ILECOMP Y����������SETUP2 Z�����  N� %��_AP2B�CK 1[� � �)��Y�h�%O������z����� N��r�ϖ��=�̿ a��ϗ�&ϻ�J��� �π�ߤ�9�K���o� �ϓ�"ߠ���X���|� �#��G���k�}�� ��0�����f����� ��,�U���y������ >���b���	��-�� Qc����:� �p�);�_ ���$�H�� ~/�7/�D/m/� �/ /�/�/V/�/z/? !?�/E?�/i?{?
?�? .?�?R?�?�?�?O�? AOSO�?wOO�O�O<O �O`O�O_�O+_�OO_��O\_�_��3�P7�� 2L�*.VR�_�_DP*�_�_AS0o)oU�PPC1oZo>DPFR6:Eo�no�o9kTΠ�o�o�oe�o
|���o0VG*.F�_aCQ	qc�O�|�A{STM �r��nt`���DPiPend�ant Pane	l�A{H�i��wW�p����BzGIFŏ���uۏ����?�BzJPGI�s��u_��.��ß:jJS͟��DP���䟡�%
JavaScript"�M�CS�z��vg�$�� %Casca�ding Sty�le Sheet�s��P
ARGN?AME.DTկ8\�p\鯧�	��*��֯�DISP*  ���pm���<������Z�	PANEL1���%�p�1�$�6��2&ό��z�7�I����3����������b��4.ߔ�����?�Q����TPEINS.XML��Ɖ�:\����Cu�stom Too�lbarB�a�PA?SSWORD��6^?FRS:\��D�� %Passw�ord Config��_����E� k_i������.���R� ��������A���� w�*��`� �+�O�s� �8�\n/� '/� /]/��//�/ �/F/�/j/�/?�/5? �/Y?�/�/�??�?B? �?�?x?O�?1OCO�? gO�?�O�O,O�OPO�O tO�O_�O?_�O8_u_ _�_(_�_�_^_�_�_ o)o�_Mo�_qo oo �o6o�oZo�o�o% �oI[�o�� D�h���3�� W��P������@�Տ �v����/�A�Џe� 􏉟�*���N��r� ܟ���=�̟a�s�� ��&���ͯ\�񯀯� ����K�گo���h��� 4�ɿX������#ϲ� G�Y��}�ϡ�0�B� ��f��ϊ���1���U� ��yߋ�߯�>����� t�	��-����c��� �����L���p������;���_�q�O���$FILE_DG�BCK 1[���X���� < �)
S�UMMARY.DyGu�!�MD:�����-�Diag� Summary�����
CONSLOG������-m���Console� logn��	T�PACCNc�%�����TP A�ccountin����FR6:I�PKDMP.ZI	P!%�
9r��	�Exceptio�nv��*.DT���-�FR:\����FR DT Files��&��MEMCHECCK�J��}/��Memory D�ata~/M� `?�)	FTP`�/�d/�/�'�mme?nt TBD?M��L >))ET?HERNET�/��<!E?�?��Eth�ernet � figura����!?DCSVRF�/�/��/O�!%�0 �verify a�ll
OO�M,�5DIFF�?�?�?܌O� %!Hdi�ff�OBG<!�0CHG01�OjO|O_AX�O9_DB*��I2_��O _�_�O6_H_�B3p�_r_�_o �_�@o�VVTRND?IAG.LSEo�_�o�o�!]a Op}e�3 Log �nosticM�T�4�)VDEVabDA�zo�o!�AVis�aDe�vice�o�kIM�Gabh�o��S�9tImagE�k�UP�`ES�o~FRS:\�����Updates OList*����p�FLEXEVEN�{?����Ap� ?UIF Ev1�`���  +�l)�
PSRBWLD'.CMُ!����,�� PS_ROBOOWEL#?����HADOW����������#Shadow Chang/����L�s�RCMERR������7��#���CFG Er�ror?ptail>ڟ ��;"��SGLIB/��(�t���!�� St�0x�ad�u��)���ZD�/���;��'�ZD�`adݯj�r�NOTI�?�,�����%Notif�ic�2j�ㆀAG ��'�<�K�I�r��� ��%Ϻ���[����� &ߵ�J���n߀�ߤ� 3���W����ߍ�"�� F�X���|����A� ��e������0���T� ��a������=����� s���,>��b�� ��'�K�o� �:�^p�� #��Y�}/$/ �H/�l/�y/�/1/ �/U/�/�/�/ ?�/D? V?�/z?	?�?�???�? c?�?�?O.O�?RO�? vO�OO�O;O�O�OqO _�O*_<_�O`_�O�_ _�_�_I_�_m_oo �_8o�_\ono�_�o!o �o�oWo�o{o�o F�oj�o��/� S�����B�T� �x����+���ҏa� �����,���P�ߏt� �����9�Ο��o�� ��(���5�^�ퟂ�� ����G�ܯk� ���� 6�ůZ�l�������� C����y�ϝ�2�D� ӿh����Ϟ�-���Q� ���χ�߫�@���M� v�ߚ�)߾���_��� ���*��N���r����$FILE_F�RSPRT  ���h�������MDON�LY 1[��_� 
 ����7� �[��D��h���� ��-���Q������� ��@R��v�) ��_��*� N�r��7� �m/�&/�3/\/ ��//�/�/E/�/i/ �/?�/4?�/X?j?�/��??�?A?�?�?��VISBCK�����*.VD�?9O�0�FR:\@ION\DATA\$O��2�0Visi�on VD fileeOs?�O�O�?�O �?_�O_=_�Oa_�O �_�_&_�_J_�_n_�_ o�_9oKoooo�_�o "o�o�oXo�o|o# �oG�ok�o�0 �������0� U��y������>�ӏ�b�������-���LU�I_CONFIG7 \��A8�� $ ���{ �叟����şן���w�|x�!�3�E�W� i�y��������ү� {����,�>�P�b��� ��������ο�w�� �(�:�L�^����ϔ� �ϸ�����s� ��$� 6�H�Z���~ߐߢߴ� ����o���� �2�D� V���z�������� k���
��.�@���Q� v���������U����� *<��`r� ���Q�� &8�\n��� �M���/"/4/ �X/j/|/�/�/�/I/ �/�/�/??0?�/T? f?x?�?�?3?�?�?�? �?OO�?>OPObOtO �O�O/O�O�O�O�O_ _�O:_L_^_p_�_�_ +_�_�_�_�_ oo�_ 6oHoZolo~o�o'o�o �o�o�o�o�o2D Vhz�#��� ���	�.�@�R�d� v��������Џ�� ���*�<�N�`�r�	� ������̟ޟ🇟� &�8�J�\�n������ ��ȯگ쯃��"�4� F�X�j���������Ŀ�ֿ�x��x�� � �$FLUI_�DATA ]����-���RESULT� 2^-�V� ��T�/wi�zard/gui�ded/step�s/Expert ύϟϱ������������/�A�O��C�ontinue �with Gj�anceOߊߜ߮��� ��������,�>�P� �-�-�o�0 ���o�/�.�6���a�psR��� �����"�4�F�X�j� |�����_Є������� ��!3EWi{�����������ripx���); M_q����� ����/%/7/I/[/ m//�/�/�/�/�/�/@�/��?������s�TimeUS/DST?�?�?�?�? �?�?�?OO/OAOX�Disablx� vO�O�O�O�O�O�O�O�__*_<_N^�{�7?)?;?M?_?q224x?�_�_oo%o 7oIo[omoo�oPObO �o�o�o�o!3E Wi{��^_p_�_8�_�_�_zonu0� 5�G�Y�k�}��������ŏ׏�X�EST� Eap�rn Stande��,�>� P�b�t���������ΟX���a� �{�������`�r�acces��������̯�ޯ���&�8�S��c�nect to� Network G�~�������ƿؿ�@��� �2�D�����!���E��!Y�o0I�ntroductionJ������� '�9�K�]�o߁ߓ�/ �����������#�5�@G�Y�k�}���? qϻ�����#�5� G�Y�k�}��������� ������1CU gy������:������5�� \n������ ��/"/4/��X/j/ |/�/�/�/�/�/�/�/ ??0?B?%�? I�?�?�?�?�?OO ,O>OPObOtO�OE/�O �O�O�O�O__(_:_ L_^_p_�_�_S?�_w? �_�? oo$o6oHoZo lo~o�o�o�o�o�o�o �_ 2DVhz �������_� �_+��_R�d�v����� ����Џ����*� <��o`�r��������� ̟ޟ���&�8�� Y��}�?�A���ȯگ ����"�4�F�X�j� |���M���Ŀֿ��� ��0�B�T�f�xϊ� I���m����ϥ��� ,�>�P�b�t߆ߘߪ� �����ߟ���(�:� L�^�p������� ����Ͽ�	�3���Z� l�~������������� �� 2��Vhz �������
 .��7��[�G� �����//*/ </N/`/r/�/C�/�/ �/�/�/??&?8?J? \?n?�??Qcu�? ��?O"O4OFOXOjO |O�O�O�O�O�O�/�O __0_B_T_f_x_�_ �_�_�_�_�_�?�?�? )o�?Poboto�o�o�o �o�o�o�o(�O L^p����� �� ��$�6��_o o{�=o����Ə؏� ��� �2�D�V�h�z� 9����ԟ���
� �.�@�R�d�v���G� ��k�ͯ������*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� ���Ͻ���F�X�j� |ߎߠ߲��������� ��0��T�f�x�� ������������� ,���M��q�3�5��� ��������(: L^p�A��� �� $6HZ l~=��a���� �/ /2/D/V/h/z/ �/�/�/�/�/��/
? ?.?@?R?d?v?�?�? �?�?�?����?'O �NO`OrO�O�O�O�O �O�O�O__&_�/J_ \_n_�_�_�_�_�_�_ �_�_o"o�?+OOOo yo;O�o�o�o�o�o�o 0BTfx7_ �������� ,�>�P�b�t�3oEoWo ioˏ�o���(�:� L�^�p���������ʟ �� ��$�6�H�Z� l�~�������Ưد�� �����ߏD�V�h�z� ������¿Կ���
� �۟@�R�d�vψϚ� �Ͼ���������*� ����o�1��ߨߺ� ��������&�8�J� \�n�-�������� �����"�4�F�X�j� |�;ߝ�_��������� 0BTfx� ������� ,>Pbt��� �������/��:/ L/^/p/�/�/�/�/�/ �/�/ ??$?�H?Z? l?~?�?�?�?�?�?�? �?O O�AO/eO'/ )O�O�O�O�O�O�O
_ _._@_R_d_v_5?�_ �_�_�_�_�_oo*o <oNo`oro1O�oUO�o �o�_�o&8J \n������_ ���"�4�F�X�j� |�������ď�o�o�o ���oB�T�f�x��� ������ҟ����� �>�P�b�t������� ��ί����Տ� ��C�m�/�������ʿ ܿ� ��$�6�H�Z� l�+��Ϣϴ������� ��� �2�D�V�h�'� 9�K�]��߁�����
� �.�@�R�d�v��� ���}�������*� <�N�`�r��������� ���ߝ߯���8J \n������ ����4FXj |������� //����c/%�/ �/�/�/�/�/�/?? ,?>?P?b?!s?�?�? �?�?�?�?OO(O:O LO^OpO//�OS/�Ow/ �O�O __$_6_H_Z_ l_~_�_�_�_�_�O�_ �_o o2oDoVohozo �o�o�o�o�O�o�O �O.@Rdv�� ��������_ <�N�`�r��������� ̏ޏ�����o5��o Y��������ȟڟ ����"�4�F�X�j� )�������į֯��� ��0�B�T�f�%��� I������������ ,�>�P�b�tφϘϪ� ��{�������(�:� L�^�p߂ߔߦ߸�w� �������ѿ6�H�Z� l�~���������� �����2�D�V�h�z� ��������������
 �����7a#�� �����* <N`����� ���//&/8/J/ \/-?Q�/u�/ �/�/?"?4?F?X?j? |?�?�?�?q�?�?�? OO0OBOTOfOxO�O �O�O�O/�/�/_�/ ,_>_P_b_t_�_�_�_ �_�_�_�_o�?(o:o Lo^opo�o�o�o�o�o �o�o �O�O�OW _~������ �� �2�D�V�og� ������ԏ���
� �.�@�R�d�#��G ��kП�����*� <�N�`�r��������� ˟ޯ���&�8�J� \�n���������u�׿ ������"�4�F�X�j� |ώϠϲ��������� �˯0�B�T�f�xߊ� �߮����������ǿ )��M������ ����������(�:� L�^�߂��������� ���� $6HZ �{=��u��� � 2DVhz ���o����
/ /./@/R/d/v/�/�/ �/k���/?�*? <?N?`?r?�?�?�?�? �?�?�?O�&O8OJO \OnO�O�O�O�O�O�O �O�O�/?�/+_U_? |_�_�_�_�_�_�_�_ oo0oBoToOxo�o �o�o�o�o�o�o ,>P_!_3_E_� i_�����(�:� L�^�p�������eoʏ ܏� ��$�6�H�Z� l�~�������s�� ��� �2�D�V�h�z� ������¯ԯ����� �.�@�R�d�v����� ����п����şן �K��rτϖϨϺ� ��������&�8�J� 	�[߀ߒߤ߶����� �����"�4�F�X�� y�;ϝ�_��������� ��0�B�T�f�x��� ������������ ,>Pbt��� i�������(: L^p����� �� /��$/6/H/Z/ l/~/�/�/�/�/�/�/ �/�?�A??z? �?�?�?�?�?�?�?
O O.O@ORO/vO�O�O �O�O�O�O�O__*_ <_N_?o_1?�_�_iO �_�_�_oo&o8oJo \ono�o�o�ocO�o�o �o�o"4FXj |��__�_�_�� �_�0�B�T�f�x��� ������ҏ����o� ,�>�P�b�t������� ��Ο������ I��p���������ʯ ܯ� ��$�6�H�� l�~�������ƿؿ� ��� �2�D���'� 9���]���������
� �.�@�R�d�v߈ߚ� Y�����������*� <�N�`�r����g� yϋ�����&�8�J� \�n������������� ����"4FXj |������� ������?�fx� ������// ,/>/��O/t/�/�/�/ �/�/�/�/??(?:? L?m?/�?S�?�? �?�? OO$O6OHOZO lO~O�O�O�?�O�O�O �O_ _2_D_V_h_z_ �_�_]?�_�?�_�?
o o.o@oRodovo�o�o �o�o�o�o�o�O* <N`r���� ����_��_5��_ �n���������ȏڏ ����"�4�F�j� |�������ğ֟��� ��0�B��c�%��� ��]���ү����� ,�>�P�b�t�����W� ��ο����(�:� L�^�pςϔ�S���w� ���ϭ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ������������� ���=���d�v����� ����������* <��`r���� ���&8�� 	��-��Q���� ��/"/4/F/X/j/ |/�/M�/�/�/�/�/ ??0?B?T?f?x?�? �?[m�?�OO ,O>OPObOtO�O�O�O �O�O�O�/__(_:_ L_^_p_�_�_�_�_�_ �_�_�?�?�?3o�?Zo lo~o�o�o�o�o�o�o �o 2�OChz �������
� �.�@��_a�#o��Go ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n�����Q���u�ׯ �����"�4�F�X�j� |�������Ŀֿ迧� ��0�B�T�f�xϊ� �Ϯ������ϣ��ǯ )����b�t߆ߘߪ� ����������(�:� ��^�p������� ���� ��$�6���W� �{���Q�������� �� 2DVhz �K�����
 .@Rdv�G� ��k�����//*/ </N/`/r/�/�/�/�/ �/�/�??&?8?J? \?n?�?�?�?�?�?�? ���O1O�XOjO |O�O�O�O�O�O�O�O __0_�/T_f_x_�_ �_�_�_�_�_�_oo ,o�?�?O!O�oEO�o �o�o�o�o(: L^p�A_��� �� ��$�6�H�Z� l�~���OoaosoՏ�o ��� �2�D�V�h�z� ������ԟ���
� �.�@�R�d�v����� ����Я⯡���ŏ'� �N�`�r��������� ̿޿���&��7� \�nπϒϤ϶����� �����"�4��U�� y�;��߲��������� ��0�B�T�f�x�� �߮����������� ,�>�P�b�t���Eߧ� i�������(: L^p����� ��� $6HZ l~������� ���/���V/h/z/ �/�/�/�/�/�/�/
? ?.?�R?d?v?�?�? �?�?�?�?�?OO*O �KO/oO�OE?�O�O �O�O�O__&_8_J_ \_n_�_??�_�_�_�_ �_�_o"o4oFoXojo |o;O�O_O�o�o�O�o 0BTfx� �����_��� ,�>�P�b�t������� ��Ώ�o�o�o��%��o L�^�p���������ʟ ܟ� ��$��H�Z� l�~�������Ưد� ��� �ߏ���w� 9�����¿Կ���
� �.�@�R�d�v�5��� �Ͼ���������*� <�N�`�r߄�C�U�g� �ߋ�����&�8�J� \�n�������� �����"�4�F�X�j� |������������ߧ� ����BTfx� ������ ��+Pbt��� ����//(/�� I/m//�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�/�?�?�?�?�? �?O O2ODOVOhOzO 9/�O]/�O�/�O�O
_ _._@_R_d_v_�_�_ �_�_�_�?�_oo*o <oNo`oro�o�o�o�o �o�O�o�O�O�oJ \n������ ���"��_F�X�j� |�������ď֏��� ���o?�c�u�9� ������ҟ����� ,�>�P�b�t�3����� ��ί����(�:� L�^�p�/�y�S���ǿ ��� ��$�6�H�Z� l�~ϐϢϴ��υ��� ��� �2�D�V�h�z� �ߞ߰��߁�˿���� �ۿ@�R�d�v��� ������������� <�N�`�r��������� ������������ 	�k-����� ��"4FXj )�������� //0/B/T/f/x/7 I[�/�/�/?? ,?>?P?b?t?�?�?�? �?{�?�?OO(O:O LO^OpO�O�O�O�O�O �/�/�/_�/6_H_Z_ l_~_�_�_�_�_�_�_ �_o�?oDoVohozo �o�o�o�o�o�o�o
 �O=�Oa#_�� �������*� <�N�`�r�������� ̏ޏ����&�8�J� \�n�-��Q��uڟ ����"�4�F�X�j� |�������į����� ��0�B�T�f�x��� �������ΰ��ǟ ɿ>�P�b�tφϘϪ� ����������կ:� L�^�p߂ߔߦ߸��� ���� ��ѿ3���W� i�-ߐ��������� ��� �2�D�V�h�'� ��������������
 .@Rd#�m�G� ��}���* <N`r���� y���//&/8/J/ \/n/�/�/�/�/u� ��/?�4?F?X?j? |?�?�?�?�?�?�?�? O�0OBOTOfOxO�O �O�O�O�O�O�O_�/ �/�/�/__!?�_�_�_ �_�_�_�_oo(o:o Lo^oO�o�o�o�o�o �o�o $6HZ l+_=_O_�s_�� �� �2�D�V�h�z� ������ooԏ���
� �.�@�R�d�v����� ����}����*� <�N�`�r��������� ̯ޯ�����8�J� \�n���������ȿڿ ����ϟ1��U�� |ώϠϲ��������� ��0�B�T�f�wϊ� �߮����������� ,�>�P�b�!σ�Eϧ� i���������(�:� L�^�p���������w� ���� $6HZ l~���s���� ���2DVhz �������
/ ��./@/R/d/v/�/�/ �/�/�/�/�/?�'? �K?]?!/�?�?�?�? �?�?�?OO&O8OJO \O/�O�O�O�O�O�O �O�O_"_4_F_X_? a?;?�_�_q?�_�_�_ oo0oBoTofoxo�o �o�omO�o�o�o ,>Pbt��� i_�_�_���_(�:� L�^�p���������ʏ ܏� ��o$�6�H�Z� l�~�������Ɵ؟� ������S��z� ������¯ԯ���
� �.�@�R��v����� ����п�����*� <�N�`��1�C���g� ��������&�8�J� \�n߀ߒߤ�c����� �����"�4�F�X�j� |����qσϕ��� ���0�B�T�f�x��� �������������� ,>Pbt��� ������%�� I�p����� �� //$/6/H/Z/ k~/�/�/�/�/�/�/ �/? ?2?D?V?w? 9�?]�?�?�?�?
O O.O@OROdOvO�O�O �Ok/�O�O�O__*_ <_N_`_r_�_�_�_g? �_�?�_�?�_&o8oJo \ono�o�o�o�o�o�o �o�o�O"4FXj |������� �_��_?�Q�x��� ������ҏ����� ,�>�P�t������� ��Ο�����(�:� L��U�/�y���e�ʯ ܯ� ��$�6�H�Z� l�~�����a�ƿؿ� ��� �2�D�V�h�z� �Ϟ�]��������Ϸ� �.�@�R�d�v߈ߚ� �߾������߳��*� <�N�`�r����� �������������G� 	�n������������� ����"4F�j |������� 0BT�%�7� �[�����// ,/>/P/b/t/�/�/W �/�/�/�/??(?:? L?^?p?�?�?�?ew ��?�O$O6OHOZO lO~O�O�O�O�O�O�O �/�O _2_D_V_h_z_ �_�_�_�_�_�_�_�?�o�?=oKi�$FM�R2_GRP 1�_Ke� ��C4  B]�P	 P�o��l�`F@ �eE����b�a�Z�a�L��FZ!D�`��D�� BT���@����m?��  �\�`6����)r��5�Z�f5�ES9q�mAg�  Qc{BHKt��`}q@�33@��p�s�\�d��}�`@�q��n�
��a�<�z�<�ڔ�=7�<�
;�;�*�<����m8ۧ�9k'�V8��8����7ג	8(���r��o�����̏���W_b_CFG `lkT�b,�>��P�b��NO ^lj
F0�� ����RM_CHKTYP  \aPt`�v`,`^aROM��_�MIN��S������pX_`SSB��aKe �f�U�0�B���TP_DEF__OW  Ttc>W�IRCOM��h���$GENOVR/D_DOؖQ���THRؖ d��dޛ�_ENB�� ^��RAVCecb��� ��eH�3���W��le�v��z [���OUh`hll����hl��e<������5�>SC�  D^�d��׶Ϗ�@�av�B���a|iعI���SM�Teci	�x`�Z���$HOSTC�19jli��_�`� MCTr��0�V  27.�0��1i�  e `߭߿������ڛ���&�8�J�m����	a�nonymous@q��������� /��`����^�`�M��� q��������� ����� 6���~�[m ����8� ��4 V�EWi{��� ����
@R// A/S/e/w/���� ��/*??+?=?O? �s?�?�?�?�?�// �?OO'O9OKO�/�/ �/�O�?�O�/�O�O�O _X?5_G_Y_k_}_�O "_�?�_�_�_�_oTO fOxO�O�_yo�O�o�o �o�o�o,_	-? Qto�_�_���� �(o:oLo)�`M��o q�������nd�ݏ� ��6�7�~[�m�� ������� �"��� V�3�E�W�i�{��� ��ïկ�
�@�R�/��A�S�e�w����EN�T 1k�� P�! ���  �� ���ؿ�п1���U� �a�<ϊϯ�r��ϖ� �Ϻ����?���u� 8ߙ�\߽߀��ߤ߶� ���;���_�"��F� |���������%� ��1��Z��B���f� ������������E�i,�P
QUICC0�v����1���9�2�:(�!ROUTER�fx�!PCJOG���!192.�168.0.10���CAMPRT,*//!%1# Q/8&RT�U/g/�/��NAME !��?!ROBOC/�/�S_CFG 1j��� ��Auto-sta�rtedєFTPܟa1����?)� �?�?�?�?�?��O.O @OROu?cO	O�O�O�O �O�O��:?L?^?;_rO �?R_�_�_�_�_�O�_ �_oo%oH_�_[omo o�o�o�o��̟ޟ� 4o!h_EWi{� To������ /�A�S�e�w����o�o �oя���<�+�=� O��s���������ޏ `�ڟ��'�9�K��� ����ȏʟ����ۯ� ���#��G�Y�k�}� ����4�ſ׿���� �f�x���gϞ���ү �������Ϭ����-� ?�Q�t�u�ߙ߽߫� ����(�:�L�^�`�2� ��q�������� ����%�H���[�m� ���������� ��� 4�!h�EWi{� T�����
��/ASew?� _?ERR l�*���PDUSIZ � ^6 ���>�WRD ?�(5���  ?guest/�/+/=/O/a/�$SC�D_GROUP [3m(< ,1"wIFT�.$PA�.wOMP�. �.�_SH�.ED�/ �$C�.COM�T�TP_AUTH �1n� <!iPendanm'�x>#;-Q!K?AREL:*x?�?�=KC�?�?�?�0�VISION �SET� (O�?,V! ?O-OWO�3{OiO�O�O��O�O�O_�O�NG4C�TRL o��aX
qQFF�F9E3_��F�RS:DEFAU�LT�\FAN�UC Web Server�ZtQ� J1�$/\�_
oo.o�@oRo�WR_CONFIG p�%��c�_�I�DL_CPU_P5C�PB����`w BH�eMIN�l��!�eGNR_IO����`NPT_SIM_DO�f�{STAL_S�CRN�f �zT�PMODNTOL8<w{�QRTYx�a�	v@K0ENB<w��#�cOLNK 1q�� ������&�8��rMAST�E�`�y`R�qSL�AVE r�H� D�uSRAMC�ACHEV�h�M1O�_CFG���s��U�O'@����CMT_�OP�P�b��YC�L��ʅ�P_ASG� 1s�g�
  :�]�o���������ɟ ۟����#�5�G�B��0�NUM��
欂IP����RTR�Y_CN��ʅ8q_�UP����q�� ج�׀��tT_  �0aT��`RCA_ACC 2u�+�  L[T� � ۪ 6P 4�� 6�-qT:�5K�  �`J�<���k���BUF001 2�v�+= 0u^�u0<��K��UV��d��p��|��߀ � ������&�3�A��N�Z�h�t�����=� �JE�UE�cu�0�r`��Z_�p��EĖE�U�EįEĻE��E��Խ�So2��2��S��Ĕu0!��SpS�u0X�]�S���ȥ���u0�p�S����T�q  �WqT ��/��@���d�  �T�z�ċ�Č�`[�~4�~u-Ԅ-�U�-Ԝ-ԫ-Ը-�U�-��-��-��-�U�������$����2������ñ��̰ ��԰��ܰ������ ������������� ��������$���,� ��4���<���D���K�<M�S�``�[�P� d�P���s�P�|�P�� P��P��P��P��𽱫�����e  ������������������������������W��������<��U (��� $�%�+ѽ�3�8�<�8� D�8�L�8�T�8�\�8� d�8�l�8�t�8�|�8� ���Ҍ��Ҕ��Ҝн���3�߹��� r̲��  rܲ�� r���Br�� 
�Br��Br�*�Br ,�:�Br<�J�K�Z� Y\�j�Y��sÂ�Y ��Y�¢�Y�²� ��²�������� ������������ ����
������ *��!+�:�9<�J�9 L�Z�9\�j�9l�z� 9|Ҋ� r�Қ� r������2w�+ 4�a\lU�!� <� p���b�HIS���y�+ �:� �2018-02-27�&�S/e/w/<�'<� : �r�/�/�/�/�/�'LN��,'1�;/(?:?L?Ѓ��'B�X�!; � `a4hq4pa4x�a4�q4��r3���cP9��?�? LM��8�W?
OO�"C<��<O�"x2:~?��2�1a4�a4�a4�ha4��a4��6O. 2L��82�?�O �O_�Yh2Y@p2�x:���2u0�:yO�Oa4��ڦO 2K�81��O�_�_�_\>u0S!0r3oo�!�oGoYo�&J�n8��_��o�o�o`2Y@�U(]f��_�%�BY@��nVC�.I�0,'09�oq���JL5_�>XZu0���o�]� 
&��/(/bp�������<�:�c��ҏ� ����/?c�P�b��oB�dh0��p09adx0 ��\@���0���0���0 ���0���0=qds�� �?�?A�.�@�.F��G� NFВ������XP��`P ��hP�������@���@ \��O�O��%�]В p0�������0������ �����P̯�_�_ݿ� π���`���B�0d ,�m��moo������ �YВ!�M��`��)�;� )wВ8pПM_�ߧ�(����IK;��b]��� }����p�5�#�5��� ;�M��ߕ����� ������)�;�)� ��q�����^4U� p2 QE� \B� �� �0 �0����0���
 ��
�e�Rd-I�KK ���"�2��"XR� `R � hR� pR-u� �B� �;(:L]��� ���S���/ /(/��cR/d/-i�/ �/�/�Ϧ��/�/ ?7/ m<��b>?P?b?�
8r �?t��/�?�?�?�?������rJO\OJ�I_CFG 2za�� H
Cycle Time<��Busy:��Idl�B�Dm�i�<�AUp|�F�ARead�G�Dow�8�O ��B�CCoun}t�A	Num �B"�C�dKF]<�Q,��SDT_ISOL�C  a�� ��PgNJ23_DS�P_ENB  �}Ze�POBPRO�C�S�E�S�SOG�_GROUP 1�{}[��< �GP?.E<�odOE?:�W_Jo<�Q`o �o�o�oho�o�o�o�:��_�X�PIN_�AUTO�T�W�SP�OSRE�_�VKA�NJI_MASK�ivQzKARELMON |a�O_<�y�o����)�gN�r~B}a���R�A<�K�fxuCwL_LApNUM�P���}pEYLOGOGING}�f������UmPLANGUA_GE a����DEFAUgLT ��O�LGA�~Y��s �~���  8�@*���<�'GI�<���9��B<�;��
�c�(UT1:\9��� �������� ͟ڟ����"�4�]��(���J�LN_D?ISP }[�L�_o]o��OCTOLL֠<�DzgP�QA���OGBOOK ��(�W��AW�W�(�rV�H�Z�l�~����������CĹ��	�
�Q�a�F���E��_BUFF 2=�}[ �S�'�i�o��G�ϝ� ������ ���	�6�-� ?�l�c�u߇ߙ��߽�����߮�7�DCS ����R=��� �� �_�Ed�v����IO 2��C �@��@gP��� ������+�=�O�c� s��������������� ';K]o�~��ER_ITMz^d!�� $6 HZl~���� ���/ /2/D/�N�SEV}����TYPz^��/�/8�/S-bqRST����SCRN_FL 32���0�D�D?�V?h?z?�?�?�?�/T�P��z_�"�NG�NAM�T�E��U�PS��GI� ���UA_LOAD��PG %�:%;DFC@GI6�?�[�MAXUALRMX����@��U
�BN%A_PR*D� ��4Q�@C�����O�t�wM�@�PP 2�.� �"f	�/I_ 4_m_X_�_�_�_�_�_ �_�_�_!ooEo0oio {o^o�o�o�o�o�o�o �oAS6wb �~������ +��O�:�s�V�h��� ��͏�����'�� K�.�@���l�����ɟ ۟�����#���Y� D�}�h�������ׯ¯ ��ޯ�1��U�@�y����n�����ӿ|HDBGDEF ��5�8��O�_LDXD�ISA
@�;��ME�MO_AP@E {?�;
 � ��]�oρϓϥϷ�����τ@ISC 1�
�9�@�ƿ(�´π>���w�bߛ�
���_MSTR �l-~��SCD 1�L������1��U�@� y�d�v�������� ����+�Q�<�u�`� �������������� ;&_J�n� �����% I4Fj��� ����!//E/0/ i/T/�/x/�/�/�/�/ �/?�//??S?>?c? �?t?�?�?�?�?�?�?�O��MKCFG ���ݗ@XO�@LT�ARM_@B�WVB*PB���O�D�@�METPU(�Bۆ���NDPAD�COL�E��NCM�NT�O �EFNp�@�O�G�� ����K^�C�Ac_mT�EPO�SCFW^PR�PM�O}YST�@1���� 4@@<#�
�QA�U�_g �_ooo[o=oOo�o so�o�o�o�o�o�o�o�3'iSq�ASI�NG_CHK  �_$MODAQ�sC��TKVN�uDE�V 	��	M�C:�|HSIZE�(�@ȣuTASK� %��%$12�3456789 �D�V��wTRIG �1��� l��% �̡�C��ˏ����&��YP����t�sE�M_INF 1��zG�`)AT&FV0E0؏�O�)7�E0V1�&A3&B1&D�2&S0&C1S�0=>�)ATZO�����H��ϟ^�Ï����A��'��K�2�o��� 5���Y�k�}� �� ���$�[�H�Z�� ~�9�������ؿ���� ���ӯ�V�a���� ÿ��k�u��ϡ�
��� .�@��d��)�;�M� ��q���������<� ��`�r�Y��I�[��� ߑߣ��&���J��� n�)�3��_������� ����"�������| /�����������0T�NIT�OR4PG ?�{ �  	EXESC1C�2�3�E4�5�g��7�8�9C�$ �$�$�$�$ �$�$�$�$T�#2	(2(2!(U2-(29(2E(2Q(U2](2i(2u(3	(�3(3��qR_G�RP_SV 1��$� ([q���>�X�<��ڴ0+&��C��?���}.�_�D��]3ION_�DBB@��}A � �@�x�5ƫ;�@V�A  �N B�?�y-ud1�uO%O7OjA�PL_NAME �!;U`@�!�Default �Personal�ity (fro�m FD)�1�AR�R21 1�L?68L@P`A�0
 d^R�O�O�O �O�O__+_=_O_a_ s_�_�_�_�_�_�_�_oo'o�s2�ORodo vo�o�o�o�o�o�o�o�r<Ao0BTf x������?H$BAB�
�B�ADP1�n��������� ȏڏ����"�4�F� X�j�|�K�]���ğ֟ �����0�B�T�f� x��������������� ��,�>�P�b�t��� ������ο����� H�6 H?�b H\�AG70"�0�C�U�ABd?�'� tφ�jϨ϶�(��=J���������!�$� �<�2�D�V�t�z߀�ߺ�70�����AB�	`&� �2�D��:�oA�Bd�v����� A� � ��B�C�XI�0��@ � �J`@�� @D� M ��?�����?A@���AAA��6Ez�  ��~?H;�	�l�	 ��@� c020�0E� ����� � � ��j�70J��K� ��J˷�J�� �J�4�JR�<ܚ5�T����70@�S�@�;�fA6A���A1UA���X�����=�N���f������T;f��X���ڤ��*  ���  �5��>6 ���5Ȭ�N0��?���#��AA����5� ����������ҍ z0� (*�0�� �0����
��	'� �� (I� ��  ����:��ÈLÈ=����d���� �<E�� �� � � ���=K����8u�1�  '�0$��� @!�p@�Wa�@ @ @![C5 CF �F �A B��CI�1��@����������A�����_�_��@A@�%AAD���/�/? ?>?)=u�i!y5AC�� :��  >�x?�ff�Ϫ?�?N? ���?K���8A@O'J>�� ���� TFP^Hy9�[�T�T��>�����1�<2�!<"�7�<L��<`�N<D��<���,���O�?������DB��?fff?�� ?&P��@T���Q?�`?U?ȩ?X�(Q� p"Q�P
��\_��{_ �G@��?�_�_�_�_�_ �_oo@oRo=ovo�EUF� eo�oao�o�M_�oqY�o*�hHm�N H[��G�� F��3l~ i������� ��D�/��m�1�� �o��ڏM����"� 4��OI�[�����y�����֟���"q  ���� CП5�̟Y�D��\ �c�j�������e����q�BHF E�R ��P��}��|� �@Iܸ�@�n�@��@�: @l��?�٧]� ���%�n�������=�=D���T�f���@��oA�&{C/� @�U|��
 +J8��
H���>��=3H���_�� F��6�G��E��A5F�ĮE���̿ް��f�G��E��+�E��EX����ް>\�G�Z�E�M�F�lD�
����i� Tύ�xϱϜ������� ����/��S�>�w�b� �߆߫��߼������ �=�(�a�L�^��� �����������9� $�]�H���l������� ��������#G2 kV{����� ��1.gR �v�����	/ �-//Q/</u/`/�/Є/�/�/��(��43��/�A��5�%�3�ϩ�/?�4� �{ ?2?��0�+#L?^?@2jb�x?�?1E�䴛|�@�;�9�?�?O�?(,OL��P�BP^Nm�z��O�/�O�O�O�O�I�0��O�O'__7_]_H_�$`_r_�_�_ �_�_�_�Ol�&ooJo8lePoZo�o~o�o�o�o�a)�o�o�8&\jz  2 oH�6�H��2�s\��B	���ݠSB���A�@� ��֣���'�9�����y�������T���Tt����Q�xv�
 ɏ�+�=�O�a�s� ��������͟ߟ��܂�� ��H;����4�$MR_C�OM �HH���z�3yG%�% 234567O8901c�u� `�H�����0�0ݡ�0��1
����not sentc *먒1��WPE�TESTFE�CSALGRm`gD�:�qd(�灿�
8�kp�t@�4#�U��S�e�w��� 9U�D1:\main�tenances�.xml��ؿ  ����DEF�AULTA�<�GR�P 2�G� ��p~�5  �%�1st mech�anical c�heck���1�Ft��|Å�lu;@ H����������ϒ2L��controll�er\�&�u�J�mt���v߈ߚ߬߾���MS��ߒ2"8���0��lue�2�D�V�h�z���C߬������)����"�4��F��CU�geQ�.� batteryJ����lu	�����������
�Sup�ply grea�soa1�3��H<�0RYlu����Ъ���^�caCbl.E���
u J\n��Y��i���9/ /2/ D/V/�Q�~/�<LH�/ �B��/�/�/	??j/ ??�/�/�/s?�?�?�? �?�?0?OT?f?x?MO _OqO�O�O�?�O�OO �O>O_%_7_I_[_�O _�_�O�__�_�_�_ o!op_Eo�_�_{o�_ �o�o�o�o�o6oZo loA�oew��� �o� 2�V+�=� O�a�s������͏ ����'�9���]� ����Џ⏷�ɟ۟� ��N�#�r�����W�}� ������ů��8�J� \�1�C�U�g�y�ȯ�� ������"���	��-� ?ώ�c�u�Ŀ��追� �������T�)�xϊ� _߮σߕߧ߹���� ��>�P�%�t�I�[�m� ���ߵ�����:� �!�3�E�W���{��� ��� ������� l�A���������� ���2Vhz ;as����� .@/'/9/K/]/ �n/�/��//�/�/ �/?#?r/G?Y?�/}? �/�?�?�?�?�?8?O \?n?CO�?gOyO�O�O8�O$K�2	 @�O�O �O&O_._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o��o�o�o�o�o � �\A?� �C _=Oa�6)p����8*�** 6A8F}p���*��N�`�r�����_OXC���Տ� �����/�A������� �������	�˟��� �c�u�۟a�s���ϟ Y���ͯ߯)�;�M�� 9�K�]������������6�$MR_H�IST 2�4E���� 
 \B$� 2345678�901��ֿ�r�9�?k�}�4�f��? �����Ϡϲ��1�C� ���Zߋߝ�T���x� ���߮����?�Q�� u�,���b������ ���)���M�_������SKCFMAPw  4E��U~r;�;������ONREL  �;�������EX_CFENB��
�����FNC��JOGOVLIM��qd��O ��KEY���R[_PANp��mi��RUNB�nSFSPDT�YP&����SIG�N����T1MOT�D����_CE_�GRP 1�4E����@P;�= z�d�\��� ��/5/�Y//R/ �/F/�/�/�/�/�/? ??C?�/M?y?`?�?�T?�?�?�?�?�;��Q?Z_EDIT�����TCOM_CF/G 1���	VO�hOzO 
7A_AR�C_�1	T_MN_MODE���	UAP_C�PL�ONOCH�ECK ?�� �� _&_8_ J_\_n_�_�_�_�_�_��_�_�_o"o��NO_WAIT_L�l,GNT?A�����5;�ta_ERR&!2�����|�o �o�op|��&Oe�@�O�c��m|  ����183��A���?�0,8��]�·��B����9�<� v� ?��7��,��n�bP�ARAM�b����v�?��w��1�C� = G�`�r�z� T������������ҏ0�,���w�^�p������CUM_RSPACE����}A͟�ה�$ODRDS�P�C�OFFS?ET_CAR"@�O�
�DIS��S_�A�@ARK�-IO�PEN_FILE�6��}A-F�PTION_IOcu���M_PRG %���%$*ǯٮj�WmOV��'s�v�
�;�t�  ���u$���$�	 a�9�$��;����RG_DSBL  �����j���RIENTTO���;�C����A ��UT_SIM_ED����r�V�?LCT �~m)B��՝;�Z �_PEqX�@9�(�RAT�G� d(��UP� ��}������Ϝς������$P�ALxb�~n��_POS_CHW�5�����p2 �L68�L@Pݳ
 d��R�d�v߈ߚ� �߾���������*� <�N�`�r�����9�2A������ �2� D�V�h�z����s��� ��������"4F Xj|�>�aǓ�y�����bP� *<N`r��� ����//�� J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? '/9/�?�?�?�?�?�? �?OO0OBOTOfOxO`�O�O�}?�w��O�M"Â�_^_@_ NW�M�M���_|_�_hW%��W�_�_�_�_o o0oRo�P��uo�l
t�T	`�_�o�o�o�a:�o±�o|0�PA�  Gy��'�Op�1������� 6�>�b@ �^���~}p @D�  �q��q�q|q?� �q�D�  Ez�s���;�	l�r	 ��@� 0@�A��p� ��p� � �� ���PH�0#H��G���9G�ģG�	{Gkf�àWT���OP�b��PCᷰ���p&�D	� D�@ D�w?������  �5��	>���pú�������� B��Bp{��!���O	ߔ��R �&��q;�0�S�K��\�)���p�(  �
p���Ј��_���U	'� � Ē�I� �  ��Hp�[=����������� �<�p� �� � � `�_�:��_�D�k�r�Nð��  '԰h��u��C��C���݀B�p������ʯ� ސ��@�2�����.�����G}±�nDp@� h��r�u����}� ����ڿŽ�#��Ş�� :��>8�x?�ff__F�X�� �`�ϟ�ѱ�8� ����>�� 8��qȺ���P�����q�s�tZ�>����<�@�<2�!<"�7�<L��<`�N<D��<���,(�e�tϖs��N���Dp?fff?�h�?&��ʹ@T�����?�`?U?ȩ?X��Ѽ	 ��ѩtȹ�u�ߖw� ���tw�L�7�p�[�� ����������$� ��H�3�l�����e����a�HmN H[���G� F����>)b M�q����� o�	�[���O��v �����o�����*//N/9/r/]/`P���"Ht�/ Cl/��/h/�/�-?��`�/???*?��ç�s�©-��H����O?<4�01�1@�I���@n��@��@: �@l��?٧]��? ��%��n�߱���=�=D���?�@��@�o�A�&{C/� �@�UO ��+J8��
H���>��=3H���_@O F��6�G��E��A5F�ĮE���hOz@��fG���E��+E��EX��O�z@>\�G�Z�E�M�F�lD�
�p�O�?_�O )__M_8_q_\_�_�_ �_�_�_�_�_o�_7o "oGomoXo�o|o�o�o �o�o�o�o�o3W B{f����� ����A�,�e�P� b����������Ώ� ��=�(�a�L���p� ����͟��ʟ��'� �K�6�o�Z������ ɯ���د���5� ��2�k�&B((A4��o�(�����X�3��ϩ����A4 ��{��οA�0+q#���ܲjb��&�1E�䴛| ��B�@ɀ�nϤϒ��ϔ��)P`�P��- #�v�/�Y�D�}�h�A���ߊ��߮�������B$���G�2�k� V��6��������e����,��<�b�P�.)h�z������������
  2 7H�6FH�;�'�\�FB�!�!y0B)Ȏ0�0A@@�/n�������/ ��'9K]D���@@�r@E
 e �����/!/3/ E/W/i/{/�/�/J�� ������4��$PARAM_MENU ?@���  �DEFPU�LSEK	WAITTMOUT;�RCV? �SHELL_WR�K.$CUR_S�TYL0B<OsPTXX?PTBm?�g2C=?R_DECSN0�ž<�?�?�? O OO$OMOHOZOlO��O�O�O�O�O�!SS�REL_ID  �<����EUSE�_PROG %��*%�O>_�CCCR�0�B��#QW_HO�ST !�*!VT�_KZT�]_�Sv_�Q�S�_J[_TI�ME2�FfU� GDEBUG�@�+�C�GINP_FLM3SKoCiTRRoCgWPGAp` 3l��kCHQoBhTYPE�,� �O�O 1,>Pyt�� ����	���(� Q�L�^�p��������� �܏� �)�$�6�H��q�l�~�����EeWO�RD ?	�+
 �	RSq`���PNS��Q4��J9O�1��TE�P��COL�յ�@��g�TRACECTL� 1�@��!+ ���������d�DT Q�@�����D � ��ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/� A�S�e�wωϛϭϿ� ��������+�=�O� a�s߅ߗߩ߻����� ����'�9�K�]�o� ������������� �#�5�G�Y�k�}��� ������������ 1CUgy��� ����ï#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/Se w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q�G�� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�3��$PGTRACELEN  �1�  ����0��6_UP �����A�
@�1@�1_C�FG �ET�3�1@�/D/D�IOTG�0TJ  ��TEBDEFSP/D �"L�1�0���0IN@TROL �"MBA8cE��APE_CONF�I@�E��A/DTI�0LI�DC�"M	XGR�P 1��G� l�1@� � �[��1A?�x�D P�D�V�C2��WO��0dcD�Y�Y�A�@�&PTOeBfK�_G ´�S�_�[B�P a�_�_�_$ooHo�1�>'oY>a���fo�o�n�o =N�=R�o�o�o �o%I4�oX��T���  Dz�s��0
���-� S�>�w�b��������� �Ώ����=�(�a��o�)�1
V7.10beta1/D���B(�A�\)A�G�NQޚ�>�ײ������A����ff��A��p�AaG�?�  ޑ@��OP��� o���+�=�/CA	p��^b�D�u��������CQKNOW_�M  _E*F
TS�V �9Y��E
���1�J��U�@�R���/B�]	SMR2S���0���	AE?���p����l�BD������@zA��.�6�2�XD̲�
QMR2S���TVi���_d�Ϻ��M{ST2Q1 1�I��4�E�Ȫ�� ^F��	��L�?�Q�c� �߇ߙ��߽������ �J�)�;��_�q��������2��ͱ�ώ�0�< ���3P3 
��.�@���4]�o�������5�����������6'9��7 Vhz���8�������MAD�6 �
F��OVLD � K���P�ARNUM  p�ˁ���SCHN	@C
����3%UPD��UO/>��_CMP_���0�@�0'*Eg$ER/_CHKu%(CBB�&r/�+RS��ů
QG_MOP�/�%_�/~��_RES_G���K
���_d?W?�? {?�?�?�?�?�?O�? *OONOAO4&5	�1<A?sO&5\�O�O�O (3���O�O�O(3 _ -_2_(3U M_l_q_(3 � �_�_�_(3� �_�_<�_(2V 1���1�ͱ@`|��"T?HR_INR0!���5d^fMASS6ko ZgMNjo�c�MON_QUEUE ���Φ0c�U 4Nl U�!N�f�h�cEND�a?y�EXEu1 BE�p�o�cOPTIO��g;�`PROGR�AM %�j%��`)o��bTASK�_IPb~OCFG� ��o���pD�ATA��� �@#�2صf�x����� ��Y�ҏ�����ŏ�>�P�b�t�'�INFO���D���d0�͟ ߟ���'�9�K�]� o���������ɯۯ�@���#�5������D�� _I�q� DIT� � ������tW�ERFL<xQc��R�CALL_CON�F Ƅ�����%�0�@�R��ʶݳKN�p?�� 0�ڶLDB�D 1��.��]���/���VL dp�%�7�I�[�m�� �ߣߵ����������� ��&���J�\�n��� ���A����!�� ��&�8�J�\�n��� �����������!�� ����2��Qcu� !������ ,>Pbt��� ���//�7/ I/[/��//��/�/ �/�/ ??$?6?H?Z? l?~?�?�}/�?��? �/OO/OAO�?hO�? �/�O�O�O�O�O�O
_ _._@_R_d_v_�?�_ uO�_�_O�_oo'o �_No�Oro�o�o�o�o �o�o�o&8J \7o��_��)o� ��1o"��goX�j� |�������ď֏��� ��0�c�f���� 9�����ϟ�O���� M�>�P�b�t������� ��ί����I�:� �3�p���������ǿ a��!��$�6�H�Z� l�~ϐϢϴ������� ��׿ �S�D�V�ɿw� �ߛ�ѿ��Y����
� �.�@�R�d�v��� �����߽��9�*� ��K�]�o������?� ������&8J \n������� ���C�1CUg �������� //0/B/T/f/x/�/ �/w�/��/�/i? )?;?qb?�/��?�? �?�?�?�?OO(O:O LO^OpO�/]?�O�/�O y?�O�O_!_�OH_�O �?~_�_�_�_�_�_�_ �_o o2oDoVo�Ozo U_so�o�O�o�o�o �o.a_Rdv�� �������*� <�`��o����	�� ɏۏ���G8�J� \�n���������ȟڟ ����C���F�y�j� ���������/��� -��0�B�T�f�x��� ������ҿ���)�� ���Pσ�qσϕϧ� A��������(�:� L�^�p߂ߔߦ߸��� �߷� �3�$�6��W� i�{�Ϣ�9������� ��� �2�D�V�h�z� �������ߝ����
 ��+=Oa��� �����* <N`r����� ���#/#/5/G/ �n/��/�/�/�/�/ �/�/?"?4?F?X?j? |?W/�?��?�?I/�? 	OOQ/BO�?�/xO�O �O�O�O�O�O�O__ ,_>_P_�?=O�_�?�_ YO�_�_�_oo_(o�_ mO^opo�o�o�o�o�o �o�o $6i_Z 5oS��_���� ��Ao2�D�V�h�z� ������ԏ���
� ��@�sd�v���� ������y�'��*� <�N�`�r��������� ̯ޯ�#�ݟ&�Y�J����k�}������ �џҿY���� ,�>�P�b�tφϘϪ� �������Ϳ�9�:� �[�m�ߑ��ϸ�O� ���� ��$�6�H�Z� l�~���������� ���� �S�A�S�e�w� �������������
 .@Rdv�� ������y�' 9K��r	���� ���//&/8/J/ \/n/�/�m�/��/ ��/??1?�/X?�/ ��?�?�?�?�?�?�? OO0OBOTOfO�/�O e?�O�O�/�O�O__ �O>_q?b_t_�_�_�_ �_�_�_�_oo(o:o Lo'_po�O�o�o_�o �o�o!_�oW_HZ l~������ �� �SoV��oz� )������я?����� =.�@�R�d�v����� ����П����9�*� �#�`����������� Q�ޯ���&�8�J� \�n���������ȿڿ �ǯ�C�4�FϹ�g� yϋ�����I������� ��0�B�T�f�xߊ� �߮�������)�� ��;�M�_�q��ߘ�/� ����������(�:� L�^�p����������� ���� 3�!3EW ��~������ � 2DVhz �g�����Y/ /+/aR/���/�/ �/�/�/�/�/??*? <?N?`?�M/�?��? i/�?�?�?O?8O�? }/nO�O�O�O�O�O�O �O�O_"_4_F_y?j_ EOc_�_�?�_�_�_�_ �_oQOBoTofoxo�o �o�o�o�o�o�o ,oP�_t��_� ��o��7o(�:� L�^�p���������ʏ ܏� �3�6�iZ� 	�{��������؟o� �� �2�D�V�h�z� ������¯ԯ��
� ��@�s�a�s����� 1���������*� <�N�`�rτϖϨϺ� �ϧ���#��&ߙ�G� Y�kߡ���)�׿���� �����"�4�F�X�j� |����ύ���	��� ���-�?�Q���x�� �߮��������� ,>Pbt��� �����%7 �^������� �� //$/6/H/Z/ l/G�/��/�/9�/ �/?A2?�/wh?z? �?�?�?�?�?�?�?
O O.O@Os/-?vO�/�O I?�O�O�O�O_O_�O ]?N_`_r_�_�_�_�_ �_�_�_oo&oYOJo %_Co�o�O�o�o�o�o qo�o1_"4FXj |������� ��o0�coT�f��o�� �����oҏi��� ,�>�P�b�t������� ��Ο���͏�I�:���[�m�����$P�RCALL_VE�R  ���T���WOR�K 2̰�� ?
 \G�����Q�( ��W�2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� ���� �R�0��V� |������������ ��0�B�T�f�x��� ������������ ,>Pbt��� ����(: L^p���`�� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O0���O_ �0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� &_������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������t� ʿ���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��������������س�$�PRGADJ ��ֵ�A7�  *�? 4�7��d?��NS_CF�G �ֵ��?�  Bzt?�7�@7�<@�?�k�%�k��������k�J�GRP 2��X�'� 	H W l����e��?z�A ?��t$�* / **:%7�*F ҷ`Է����?� �R�bt��� $���: Lzp����� ��h//$/R/H/Z/ �/~/�/�/�/�/@?�/ �/*? ?2?�?V?h?�? �?�?O�?�?O�?
O �O.O@OnOdOvO�O�O �O�O�O�O\___F_ <_N_�_r_�_�_�_�_ 4o�_�_oo&o�oJo \o�o�o�o�o�o�o �o�ox"4bXj�������ֶ	 :�q�\�����	 ����叀�	��H�PREF �X��7�7�
F�IOR?ITY  k�$��7���MPDSPON  ����v��UTb���K�I�OD�UCT_ID e����OG���_TGLb�!���TOENT 1�����(!AF_I�NE��2�=�!�tcp=�e�!�udT���!iccm|�����XYQ���� �?�)�a 2��7��� ,���X�?�|�c�u� ����ֿ������0�H�T�f�*��Q��X������ϻ�?�>5H�,�2/<����k������Az�,/  �N��e� w߉߭��7��?�Q��/��PORT_N�UMb�7�m���_CARTRE�P��֬H�SKST�A�� �LGS6/����z�7��Unothin�g��r���%�6�T?EMP �����-�Z�_a_seiban���� ;�&�_�J���n����� ��������%I 4mX}���� ���30i T�x����� /�///S/>/w/b/��/�/�/�/�/�/��VOERSI�&0� disab�led ?SAVE� �Ě	26�70H755�(�/�?!�τ?�?���?C 	�8��/�KOR�e$OMO_OqO�O�JA<L�?�O��F2_�W 1��o0P����u__�w0�UR?GE_ENB����lm�ǡWFKPDOb��7ү�W+�lT/���W�RUP_DELA�Y ��_UR_?HOT %T�������_}UR_NORMAL�X̒�_0o�WSEMIo5oto.�_QSKIP�Cܹ��Cx�/�o�/�o�o �m�2 Vhz@ �������� 
�@�R�d�*�t����� ��Џ⏨����<� N�`�&���r�����̟ ��ܟ��&�8�J��U�$RBTIF��	�RCVTMOU����h�DC�R�Cޗi ���a?XB����B%�>N�� @�"�ymS��`�M]y��+(��i��o� <2��!<"7�<L���<`N<D��<��K��O�x���R߮���ҿ��� ��,�>�P�b�tϤ��RDIO_TYP�E  �Mj���E�FPOS1 1�
N9��x�?��Rg�  ��D��?h�ߌ�'� ����]��߁�
��.� @�����'��s��G� ��k������*���N� ��r������C�U��� ������8��\�� Y�-�Q�u� ���XC|�ϿOS2 1�[ ��3m�i/���3 1���/��/n/�/%/S4 1�</N/`/�/??<?>�/S5 1��/�/��//?�?�?�?O?S6 1�f?x?�?�?BO�-OfO�?S7 1� �?OOYO�O�O�OyOS8 1�O�O�O��Ol_W_�__SMA_SK 1�� ��8�_�V�WXNO���V�oc��MOTE�o���T3a_CFG� �:m�Qa��P?L_RANG6ar��taOWER ���`�fSM_D�RYPRG %��Z%7_�o�eTAR�T �n�jUME_PRO�o�oI�T_EXEC_E�NB  _�z�GSPD"pdplx��{vgTDB��zRM���xI_AIRPU�R}` �_��]M�T_�PT�`8k~��h�OBOT_IS�OLC�^iffe�D�NAME ��z8��OB_O�RD_NUM ?��h�qH?755  ��֏����h�PC_TI�ME��v�xh�S2�32Sb1뮩`�L�TEACH ?PENDAN��OW�hW�6_!M�aintenance Cons���f���"��No UseW���y��ן�������2�N�PO�`�az(�/�CH_L%p3�3�R	��l�?!UD1:ǯn�=R�PVAIL�����&�.aSPAC�E1 2���k�nbO�E�USP�nb������< �@�?�﫫�﯋� ��ٿ��?�Q�c� u�'ϙ������ϑ��� ���*u.q'�C�U�g� y��ϝϿϵ��ߕ��� ���!�;�Q�c�u߇� 9����������� �;�M�_�q��5��� �����������+ I�[�m���������� ���$�EW i{�?���� � //5/Sew �;/���/��/�/ ?�/?O/a/s/�/�/ I?�/�/�?�?�??*O O?O]?o?�?�?EO�? �?�O2O�O_&_�O;_tt�&�2+�� =� sO�O�OI_�O�O�_6_@�_&oGoo\o]_3p_ �_�_�_�_jo�_o�Wo�oGh?}~o4 �o�o�o�o�o��o/ 2�x�h���`����5�������� P�S���3�����������6ӏ���	��͟ ?�q�t���T���˯����7����*�<� �`�����ۯu�˿�ÿ��8�'�9�K� ]�ρ���������������"�#�G �N9� �ZD
��7 r�  9ţ� �����������;�vȀ.�]�;�Z�ߍ�]Ad ���ߚ���������� "�4�*�<�N�?�|��� �����6���& 8J@�R�d�v���� �����V"4F Xj`r����w `� @`@�%k�/��	O!y �`/r/xR*S/�/�/ �/�/�/�/!?3?�/? ?K?�?O?a?s?�?�? �?O�?�?AOSOO'O 9OkO�OoO}
1/_�a[_MODE  �9�y�VS �"9��O����-/�V_�_�Z	�_�_�dCWORK_AD(\��
x4��aR  9�F�?`�_)`_INTVAL(P�ĐA�QfOPTI[ON`f ke�p�V_DATA_G�RP 2�D�D� P�_�o�_�o�i �O	?-cQ� u������� )��M�;�]���q��� ��ˏ���ݏ���� I�7�m�[�������� ş�ٟ���3�!�W� E�g�i�{�����կï �����-�S�A�w� e���������Ͽѿ� ��=�+�a�Oυ�s���ϻϩ���/Q�$S�AF_DO_PULS`0P�a�	���CAN_TIM'Q���e�R ����`��P{5P���҇S�a�Rg�}QY�� �o�ߣߵ��� ����z��!�3�E�W�i�sX��2H��Yѝ�d����bW�t� Cn����	��r���� �`��_ "  T�>`/�l�~�����T D���������� �� 2DVhz ������c_yU���0B��	!iў;��otzTpbe 
�t��Di�T|iђ[  � �� }Q7Qi�a�Q���� 
//./@/R/d/v/�/ �/�/�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�?�?OO&O8O�JO\OnO�O�O�Oq� ,��O�O�O__'_9_ K_]_�O��_�_�_�_ �_�_�_oo+o0am_r0*�)��|o�o �o�o�o�o�o�o 0BTfx��� ������,�>� P�b�t���������Ώ �����(�:�L��O p���������ʟܟ�  ��}_6�H�Z�l�~� ������Ư1o_eio� ��*�<�N�`�r��� ������̿ڹ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯����ߨ�������-� ?�Q�c�u����� ��������)�;�I���R�������rbx�N	12�345678��h!B!ܺ��s�|�� %7I[m� ����� &8J\n��� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??��R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO 1?�O�O�O�O�O�O_ _&_8_J_\_n_�_�_ �_�_�_�O�_�_o"o 4oFoXojo|o�o�o�o �o�o�o�o�_B Tfx����� ����,�>�P�b� t�3������Ώ��� ��(�:�L�^�p��� ������ʟ��� �� $�6�H�Z�l�~����� ��Ưد���� �q���B�T��y��������Cz  B}p��   ���}2r� } ���
���  	�q�2:�!�3�E�W�g�	��h��ϭϿ��� ������+�=�O�a� s߅ߗߩ߻������� ��'�9�K�]�o�� ������������� #�5�G�Y�k�}������h��ܲ<�� ����  ������Ƕ����t  Ѱ	 ǵ��$SCR_GR�P 1��@��#� � ��� ׵	 g�o�yi���ٵ�	���������ٰ��C����}͆$���L�R Mate 2�00iD 567�890�LRM�] 	LR2D� ds�
123	4c�v�g����oǶ^�^��D���}
��	��/'/9/K/]/Ǵ���H�o �s ^�/��/�/�/�!�s��/"?�/F?��7?j��h��,�	B���!Ƒ?�2�4�AѰ�?�  @��5�@���0�? ?�5�2H���O�:�F@ F�`2B:O1?^OIO �OmO�O�O�O�O�O _ �=�1�2+__(_:_LTB�Z_�O�_�_�_�_ �_�_�_o	oBo-ofo Qo�o|Ϛj��g�o�׷���os��1@�>��@h�0O���ew� ��9��ǴA�0�fH�u�/�%�p����s� ��$�2� ��G�S�e�4�f���
 ���������o�̏��7ECLVL  �s�����rA���*SYSTE�M*�V9.10�35 P�7/19�/2017 A� ���>�e�SE�RVENT_T �  $ $S�_NAME �!��PORT��^��ROTO���s�o_SPD{�(�� ���TRQ �  
��AXI�S������ 2��`��DETAIL�_  l $DATETI�����ERR_COD��IMP_VEL�ϰ 	�TOQ~ �ANGLES �GDISz�,���G���%$LIN�  REC�� ,肑ʕ�$�MRA~n� 2 d���IDX��i��� �f�$OVE?R_LIMI��Đ|~ ��OCCUR���  �CO_UNTER��Φ�FZN_CFG��� 4 $EN7ABL�ST ����FLAG��DEBU$�R9�(���D ��� � 
$MI�N_OVRD���$Iy�5�Y�Q�b�F�ACE��Z�SAF>y�MIXED��b��B�Y�ROB��$�NE��PP����H�ELL��	� 5$J��BAS��RSR_�  $NUM_��. � �1U���U2�3�4�5ʕ6�7�8U��R�OO��\�COy�O�NLY�`$US�E_AB���A�CKENB���I}N��T_CHK��OP_SEL_�Χ�_PU���M_v�OU��PNS�����ԳV����M�T�PFWD_KAR�����RE��$�OPTION6�$�QUE�ɝ�D�Y�Ͳ$CSTOPIg_AL��ԳEX�����j��XT��M1ڗ�2��MA^�STmY��SO��NB��;DI��TRI$�b�.�INIz�M�����NRQ�և�END���$KEYSWITCH����k��HE�BEATM�M�PERM_LE��%�E�L�U�F���S��DO_H�OMy�Oͱ��EFaP����%�АST*⚙�Ce�OM�n�O�V_MS����ET?_IOCMN��r�f����ճHK{��
 D ���S�U�`�MP���P�O��$FORC��WARN��OM��� �0$F'UNC���U����SAR��h�2g�3g�Q4\��⾠O*�LM�yw���UNLO������ED����SNPX_AS�� 0�ADD|4�6�$SIZ��$VARU�MU/LTIP����l��AM� � 1$�����	���䖒�C�IFRI	F����SJ�\���9 �NF��ODBUS_AD��	�������|� � ���6�TE��$D�UMMY8�SG�L�TA��  &����`� � �STMTj�PS3EG��BWe���SHOW��BA=NTPOFb��9�10X�����SVCy�GF� � $PC����x�£$FBI�P�S�Pr�A�����VD�zE�� �.��A00?�� p��z��������U5�6�7�8�9�A�B�[���� �F�b�(��1�1�1
)1B)1$)^��(>)1K)U1X)1e)1r)1)U1�)1�)2�2�U2�2�2
)2)U2$)21)2>)2K)U2X)2e)2r)2)U2�)2�)3�3�U3�3�3
)3)U3$)31)3>)3K)U3X)3e)3r)3)U3�)3�)4�4�U4�4�4
)4)U4$)41)4>)4K)U4X)4e)4r)4)U4�)4�)5�5�U5�5�5
)5)U5$)51)5>)5K)U5X)5e)5r)5)U5�)5�)6�6�U6�6�6
)6)U6$)61)6>)6K)U6X)6e)6r)6)U6�)6�)7�7�U7�7�7
)7)U7$)71)7>)7K)U7X)7e)7r)7)e7�)7�$ǢVPI�=U�� ��V���
R��{���o$TORS�CMX��"�M��R��ǰ �Q_ҠRx�.�ϑ%� �Φ�YSLS�|� � ����x���(��x�؄�VALAU���֨��FɁ�ID_L��9�HI�4�I;�$FILE1_��d���$��Ć�SA�� h ���VE_BLC�KMӝ����D_CPU�������g��y�ĂV���R ? � PWԠ��lp �LAS����-�&�RUN_FLG?��C�&��F�d��d�&�H��2����&���TBC2C� �� ��F������pk�Ծ���TDCF��#�עQ�b�ҧT!H�� ����R����?ESERVE��-����-�3������ X -$X�LEN��e���X���cRAIд�ȀW_����1X�Q�2��MO$����S� ��I����`]�ǹ��X�ܻDE쵞LACE�ⱃCqC��]�_MA��p�%���%�TCV,�M���T��N�m�cʯ 곖�����J����M���J�������d�2�Ћ�����*�JK�VK@������N�
�Jcl-��JJ!�JJ)�AAL�O�!�O�I�e4J�5
���N1t�P��?�)���LŰ_������CF�� =`��GROU����қN��C1��R�EQUIR��E�BUHT���$T�2�U��֞��� \��APP�R�CL��
$O�PENN�CLOSD��_�S��s��
��. �5�M�*�8�(���_MG`����C�����'���B{RK��NOLD��>2RTMO_���$���J��PQ�� !��)��m��v��%6>�7>����S�>��� ���l���!Ѭ�PATH������񄸽� r���xSCAB���O��INW�UCh˰� C�UM 	Y������'=�3��B
!�B
N�B PAYwLOA��J2LY�OR_ANߡ�L���	�}	���R_F�2LSHR'��L�O��4�4ACRL_���u(�H���$H���5FLEXQ�:��J�� P;⳯�ů,�>���RW� :d�v������y�)���������F1 �,%@'��ǿٿ����p"E�+�=�O�a� sυϗϩ�G8d4���� �T v8���������	T�7E1X��N1ճ$ �(�E�(�*�<�N� R�[�I�m�v߈ߚ߬���� ����������Z�ATY&��CEL� k�+S
�J���JE��CTR�T!TNt�'V��H�AND_VB���Q���  $�0Fi2�����SW��M�����!� $$M� �阀���X�� �\
0�U,�fA@�z ��?�#i��A�����A��A��.`��ϐ��UD��D��P��G9���iST���a���aN��DYE�L���d6e � Y�����|��4 �0�PF�O�X�@a�j�s�|����J��"�P+R���r�v���qASYM��������!0�_ ��� /���X9K]o�J�9�
p�����	f$_VI�S������V_UN!I'��>C�J�5� cu5��9��F�j�����9�,���3�BJ��H�@�a#�R�d�DI�����O
��B��C$) N@=bI �A=�4 7�Z E�E�] l���� �� % � �QME�!�@`���G�T��PT���@�������Dc������T���� $�DUMMY1N�o$PS_W RF ֊�$���FL�A��YP�3����?$GLB_T�P �����lP� XQd�&c X;��ג�ST�!��SBR��M2�1_VK2T$SV_ER� Or�^�v�SCL2�^�A� O:���GL��EW�q's 4�В�$Y�b�Z�bW������SA�a� �R��U��( ��0N۰��$G�IhP}$�� �'�P��ڰ�q) qL����q�}$Fq��E�NEAR� N�^#FKɦ TANC�^"'�JOG /� �*��$JOI�NT�1	@咤�MS�ET�q+  ��E1��!�@S�BP��@��q,� `PU��!?��LOCK�_FO� �Q�BG�LV[SGL��TE�ST_XMQ��EMP��K2�0����$U����02(�ڳ?�)
ҳP��?э'`�CE���`� �$KAR1M�T�PDRA��}�t�VcEC���x�IU?��*D�HE��TOOiL #��V$RE��'IS3���6a�T �ACH���+��O���Ҥ29ۢ��I�A�  @$RAIL_BOXE�1���ROBO�?����HOWWAR�=/����ROLM �U�A��f��A�H ��O_F�@! ����ѿq-�ΰR
��O�.�� �������OU��/�F�;�'G�1RQ��/$PIP�N�0������f ?Ѡ�CORDED���������@OG� 0 D �OBca5S���R�A�̣�A�q�7QS;YSA�ADR6Q�TCH�P 1� ,�0EN�mA
��_�����AE���VWVAc�2 Ǥ �Ч� �PR�EV_RTpq$�EDIT��VSHWR�AJ� �"��%��Dr��)>A?$HEAD����4C ����KE��Ơ�CPSPDZJM%P^�L��PR� "��3I�b��I�S6RC|PNE��7QrWOTICK #*�Mk����HN@�4� @K��Eb_GqP��nSTY����LO2�㳄��p_5 t 
��G��S%$����=J�S,@!$+��0w��4�r�P��SQUw�x%���TERC����a�PS�D6  �V��G�0�GC1��P1O����b IZ����ߡPR3��"̝��PU�A%_DYOP­�XS��K���AXI> y�D�URP�#7R6�� l��Q�P_��~�ET"P(��Z��u=F�w>A�a�Ӥ���NA��SR�T7l��YB�Z�%�V 9b�%g�#i�#/i @5Qg@5ag@5qfR5l= �iR5�<�rp9B�;~=�C�=j�|������S�SC� 8 hƃ�DS� ~�ҠSPL1�lEAT_`b !�� �ϢADDRE�S��B��SHIF��C6�_2CH6Prh�I9��A�TU9��I�Q 9��CU�STO�$AC�TV��I%�:��؀A#�p
�
���@,$NB�; \H����=\��KRC�c��"�Z��|�KQ�TXS�CREEC�<��YTINA��
��T���[��!�B�p= T�y�"~�x�U��V�L!}�L"�T��RRO�:pe�}�T �QV���UE�> ��p���9S��~�RSM� B'UNEX���Ua�S_Գuf$�eaxi�g�$��!C��Qb�T [2=�pUE�t?+�����f GMT}�L�W�[!e�O���/BBL_��W��B��@ �=rOα!rLE�B,s5��B+t�RIGH5sBRD<���ACKGR��]u�TEXn ^uYqWIDTH� U��������UI��E9Y�@qA d��z �T�!�!BAC�K��u��k�F�O*��wLAB*1?�(k�I����$UAR;����pq�Ha� B 8̑e�_B�B3�r�R������ڢ3a!�O�ApC�� ��VpUAp��R��`�LUM��c&�@'ERV��g�PO��t5Di�� GE�6�4� ��)K LPӅ�"	E�1A)��AA��QA�������5��6��7��8�����
 O�_T�Ѧ����S�C�qUSR��E �<H�q�U ��C �F�O�@ �PRI�!mx�o�ҐTRIP�m�UN�#�F���b�D%G�C%�q�6�} w G.�\��!G JTy��A�A)�OS��>�R � b���qH��³ ɾe����6�Uہq�In����cۂ �OSFF�pJF���=O�� 1H��ޤZ�I��GUx�P���!�A+��qSUB8���`SRTg��$aK�d����OR��Nq�RAU� r�T�������S��A L� HK�SHADO�W` �ӿ�_UNS�CA�ӿ��t̳DGqD�ѵ��VC"0|G��aM� �B�nF�΂���yC�� �DRIV&�!_V� Cĺ T��D~�MY_UBY }�(�De�na��Pb0���ѽ�P_հ���L%+BM(q�$� DEY��EXpp)c��t _MUx 1X(q�j`US|�� ͐�еPt��@bu�}G�0PACIN�kRG1 K�b�̣b�0��bҝc�REH��AĹѬ��bҝ�N ��@TARGh�PH�R���RU���O�p�z�M!�qQ�	�<!RmE�SWZ�_A[ђ��� O���AA(�@��"En�U0J�����p�HK5P� 3��!��Pd�sEA� n�WOR5�x���MRCV�aWQ �̀OAM5��C�S	��ޣ�ӫ�REFw����
ཀ �#�Т���������8%���Z�_RCo�[���z0Sk��t��}��dR ��p�uh���y��OU�x�� (� M��
 A2�0$�PaP � �OC A�K_ S�UL�PP��CO�I`J�Q� NT ���PE��Ob�O��O L��x��xb�̄���ĵSG� ,C�!B@ CoCACHLO������	c!�@�C�_LIMI�CFR�TX0��$HO�5���� COMM>�QbO?pG��� ρ���H@VP��i �_���ZFЏ�W�A MP�FAIjG`�� AD���IMRE��"��GPW`��� �AS�YNBUF�VR�TD6%B$�psOL��@D_ƣ^%W��PN�0ETU��� Q8��&%ECCU��VE�M~���"VIR�C�V%>#PbB!_DELA��W��鐪��AGR)R�XYZ�`c�W��3�q� T���IM�!U%�r�dT�B�qLAS�pDq�_� !��U����S �N�4E�LEXE�V�S����YA�FLZpI��(#FI` �7Ű�8��Ba����!�0��W����:�􂔊���,pORDƑ�f��C��pUX�P��T��bb��O�p���SFxp9cY  �P�O��UR粅BM�Z<����$ADJR@�3���U[��oG�2�LIN�2aXV�R�\Z2�`T_O�VR�2��ZABC^�]��3R"CwQRP��Z(��^����$�Lt��r �
�_ZMPCF^�_�B�P\d�R��LNK�rUQM�_�` ��̀Tn��TCMCM�T�C�CART_��Q-�P_|� '$J�S�TD�R�bg	�e	�/�UX!1�UUXE�@f!1e8decaIa[iIa4kf��ZZUae��JTuTZ0	�bYPD�� b.�R�ő0CHEOtРpG�W��q�0�`��c �� |D��QPWpEA�K׈�K_SHIYF��HRVFZ���<r(PCXp�R�Q! }@8�Wq�PV�Ist}D�xTRACEE��Vt��bSPHERq�d ,
 �h�o2�j�f��aFA/Z0�����|��tHOTSTA����MIPOWERFL  �� �8�WFD-O� � �q��~��1 ������/� L!��_�EIPH�����j!AFn ��ƏυO!FT������f�!��@��	��f�!R{ MAI	Ng�I��U���y�n0䂟H������!T!Pn ������d�J��!
PM�o@XYK���e9����d����f���!RDM��0V㯰�gѯ.�!OR90/���h��z�!
{�T����i�i�ƿ!RL3 C�ǿ�8���!gROS��9��4��^�!
CE�MT�Q_ϳ�kMϪ�!	"s�Cq�ϳ�l����;!s�WAS���ϲ��m��B�!s�USBC߱�n1ߎ�-� ���ߑ��� ���$�@��H��l��x�I�p�KL ?%�� �(%SVC 1�s���2���� 3����� 4�� 5�3�8� 6[�`� 7����� 8���� 9������E� ��� (����P����x�� %����M����u�� �������@���� h�����>��� f���/��0/ ���X/���/��. �/��V�/��~�/�� �x������C?�? ��?�?�?�?�?�?�? OO@ORO=OvOaO�O �O�O�O�O�O�O__ <_'_`_K_�_o_�_�_ �_�_�_o�_&ooJo 5o\o�oko�o�o�o�o �o�o"F1j U�y�������~�_DEV ����UT1�:�4��&�GRP 2��O0���bx 	� 
 ,v����O2 {�����܏ÏՏ��� 6��Z�l�S���w��� Ɵ���џ� �w�D� ��h�z�a�����¯ԯ ����߯���R�9� v�]�������п'�ſ Ͻ�*��N�`�Gτ� kϨϺϡ������� ��8��\�C�Uߒ�� ���߯��������	� F�-�j�Q������ ����������B�T� ��x�/����������� ����,P7I �m����� [��:�^E�� {�����/� 6/H///l/S/�/w/�/ �/�/�/�/ ??D? +?=?z?a?�?�?�?�? �?�?�?O.OORO9O vO�O�/�OcO�O�O�O _�O*_<_#_`_G_�_ k_}_�_�_�_�_oo �_8o�O-ono%o�oyo �o�o�o�o�o"	 F-j|c���p���J�d ��	�1��U�@�y�d������%���яQc���ꁖ����� �(��L�:�p�~��� ���f�П������ ��N���u���>��� ��̯���ޯ �V�|� M���&���n�����ȿ ���.��R�ܿF�ؿ V�|�jϠώ������ *ϴ���B�0�R�x� fߜ�����ߌ����� ��>�,�N�t�ߛ� ��d���������� :�|�a�s�*�L�&��� ��������T�9x� lZ|~��� �,P�D2h Vxz���( �/
/@/./d/R/t/ ���/ /�/�/�/? ?<?*?`?�/�?�/P? �?L?�?�?�?OO8O z?_O�?(O�O�O�O�O �O�O�O_RO7_vO _ j_X_�_|_�_�_�_�_ *_oN_�_Bo0ofoTo �oxo�o�_�o�o�o�o �o>,bP��o ��ov����� :�(�^�����N��� ��܏ʏ�� �6�x� ]���&���~�����؟ Ɵ�>�d�5�t��h� V���z�����ԯ��� :�į.���>�d�R��� v����ӿ������ *��:�`�Nτ�ƿ�� �t��������&�� 6�\ߞσ���L߶ߤ� ��������"�d�I�[� �4��|������� ��<�!�`���T�B�d� f�x����������8� ��,P>`bt ������( L:\���� ��� /�$//H/ �o/�8/�/4/�/�/ �/�/�/ ?b/G?�/? z?h?�?�?�?�?�?�? :?O^?�?RO@OvOdO �O�O�O�OO�O6O�O *__N_<_r_`_�_�O �_�_�_�_�_�_&oo Jo8ono�_�o�_^o�o �o�o�o�o"F�o m�o6����� ���`E���x� f���������Џ&�L� �\���P�>�t�b��� �������"������ &�L�:�p�^���֟�� �����ܯ� �"�H� 6�l�����ү\�ƿ�� �ؿ����Dφ�k� ��4Ϟό��ϰ����� 
�L�1�C������d� �߈߾߬���$�	�H� ��<�*�L�N�`��� ������ ����8� &�H�J�\�������� ��������4"D �������j��� ��0rW�  ������/ J//n�b/P/�/t/ �/�/�/�/"/?F/�/ :?(?^?L?�?p?�?�? �/�??�?O O6O$O ZOHO~O�?�O�OnO�O jO�O_�O2_ _V_�O }_�OF_�_�_�_�_�_ 
o�_.op_Uo�_o�o vo�o�o�o�o�oHo -lo�o`N�r� ��4�D�8� &�\�J���n����ˏ 
��������4�"�X� F�|������l�֟ğ ���
�0��T���{� ��D�����ү����� �,�n�S������t� ����ο���4��+� ��޿Lς�pϦϔ� �����0Ϻ�$��4� 6�H�~�lߢ������ ������ ��0�2�D� z�ߡ���j������� ���
�,����y��� R������������� Z�?~�r�� ����2V� J8n\~��� 
�.�"//F/4/ j/X/z/�/��//�/ �/�/??B?0?f?�/ �?�?V?x?R?�?�?�? OO>O�?eO�?.O�O �O�O�O�O�O�O_XO =_|O_p_^_�_�_�_ �_�_�_0_oT_�_Ho 6oloZo�o~o�o�_o �o,o�o D2h V��o��o|�x ��
�@�.�d���� �T������Џ�� �<�~�c���,����� ����ޟ̟��V�;� z��n�\��������� گ���ʯ�Ư4� j�X���|�����ٿ� �������0�f�T� ��̿���z������ ����,�bߤω��� R߼ߪ��������� jߐ�a��:���� ������ �B�'�f��� Z���j���~������� ���>���2 VD f�z����� 
�.R@b� ���x��/� *//N/�u/�/>/`/ :/�/�/�/?�/&?h/ M?�/?�?n?�?�?�? �?�?�?@?%Od?�?XO FO|OjO�O�O�O�OO �O<O�O0__T_B_x_ f_�_�O_�__�_o �_,ooPo>oto�_�o �_do�o`o�o�o( L�os�o<�� ��� ��$�fK� ��~�l�����Ə�� ֏��>�#�b��V�D� z�h��������� ��ԟ���R�@�v�d����ܟ�� ���$S�ERV_MAILW  
� ��樿OUTPUT����@�RoV 2��  �� (��Я\��S�AVE��TOP�10 26� d ���ο�� ��(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~ߐߢ� ����������� �2� D�V�h�z���掵YPy��FZN_CFG �����%�j���?GRP 2�燱� ,B   A�:�D;� B�;��  B4���RB21i�HELL��	����I��J������%RSR����������" F1jUg�������0_�  �>�%0�^p>|���x���uF2��d�ve�HK ;1
s� �$/ /1/C/l/g/y/�/�/ �/�/�/�/�/	??D?�??Q?c?_�OMM �s��?d�FTOV_ENB��>����HOW_REG_�UI�?�IMIO/FWDL�0�>=�^BWAIT�2���0F��6=�-IT�IM�5��gOV�A��>OA_UNI�T�3�F��LC�0T�RY�7���M�ON_ALIAS� ?e�9E�he ��"_4_F_X_fZ_�_ �_�_�_j_�_�_oo +o�_Ooaoso�o�oBo �o�o�o�o�o'9 K]n���� t���#�5��Y� k�}�����L�ŏ׏� �����1�C�U�g�� ��������ӟ~���	� �-�?��c�u����� ��V�ϯ������ ;�M�_�q�������� ˿ݿ����%�7�I� ��m�ϑϣϵ�`��� ����ߺ�3�E�W�i� {�&ߟ߱������ߒ� ��/�A�S���w�� ���X�������� ��=�O�a�s���0��� ����������'9 K]����b ���#�GY k}�:���� ��/1/C/U/ /f/ �/�/�/�/l/�/�/	? ?-?�/Q?c?u?�?�? D?�?�?�?�?O�?)O ;OMO_O
O�O�O�O�O �OvO�O__%_7_�C��$SMON_D�EFPROG �&���aQ� &*SY�STEM*>_�W� 	MWRECAL�L ?}aY (� �}/copy� mdb:*.*� virt:\t�mpback\=�>192.168�.1.103:2468 �V�_oo�)l}3x�Rfr:\�_G`�_�P�_�o�o�o9`4=eaEoWo�U�ro' }
x�yzrate 61 �o�o�o}���4e=w]}15236 ]o ��$�7{11 ���}������4e2�T:pro�g_1.tp�Uemp�^W�p���%��ݏ J�������7b9>ds:ord�erfil.da�t�_]�����,m0 �_؟P��������l��oXT�r���'� }5�oί�󯄿�� ��;M�_�q���&��9��S�P07V�032\��~ϐϢ�5�G� Q�c�u��߫���Ϗ ���ρߓߥ�8�]�\� dߩ���Ͼ����� �߅��*��N�`�r� ��'�:���K���� ������]�\�n��� #��ȟQ���v�� -�?�Z��n�#�6�=OV�7:25�44m����+n-=*.dQcl�/!/��1 ���}/�/�/4e��f\/ n/�/?#?6c1=�K/@e�/�?�?�?7b8= OZ?p0�?OO,m�_ �?�+�?O�O�O6oɿ ۹hqO__&_�o�O �Ol4u_�_�_�?�?�? ^_t_oo�_<O�_`Op�_�o�o�o }6�_|O�1052 to�o.��o�h�o }��4/F/Xj� �����/�t���� ����7�_Ro�g��� ��?oڏ�h����������$SNPX�_ASG 2����ȑ�� P 0 '�%R[1]@X栩��?���%� ��C�&�8�y�\��� ����ӯ��ȯ	��� ?�"�c�F�X���|��� Ͽ���ֿ�)��3� _�Bσ�f�xϹϜ��� ��������I�,�S� �bߣ߆ߘ��߼��� ���3��(�i�L�s� ������������ /��S�6�H���l��� ������������# O2sVh��� ����9C oR�v���� ��#///Y/</c/ �/r/�/�/�/�/�/�/ ??C?&?8?y?\?�? �?�?�?�?�?	O�?O ?O"OcOFOXO�O|O�O �O�O�O�O�O)__3_ __B_�_f_x_�_�_�_ �_�_o�_oIo,oSo obo�o�o�o�o�o�o �o3(iLs �������� /��S�6�H���l����������PARAM� ȕґ ��	�ÊP3��7�È����O�FT_KB_CF�G   �Ε��O�PIN_SIM  ț�l�~�������RVNORDY_DO  ��A���QSTP_DSBU������ـSR X�� � &�+�;�� �Y�ـTOP_ON_ERR��ׂ[��PTN X�ގ��Cx�RI?NG_PRMe�Ȓ�VCNT_GP �2W���x 	 ���֯���3���VD��RP 1��$���n��� ������ݿڿ���� "�4�F�X�j�|ϣϠ� ������������0� B�i�f�xߊߜ߮��� �������/�,�>�P� b�t��������� ����(�:�L�^�p� ��������������  $6HZ�~� ������  GDVhz��� ���/
//./@/ R/d/v/�/�/�/�/�/ �/�/??*?<?N?`? r?�?�?�?�?�?�?�? OO&O8O_O\OnO�O �O�O�O�O�O�O�O%_ "_4_F_X_j_|_�_�_ �_�_�_�_�_oo0o�BoL�PRG_CO7UNT6�玢gi'ENB��ieM�c8���o_UPD 1>�T  
Wo � �o�o72DV z������� 
��.�W�R�d�v��� ����������/� *�<�N�w�r������� ��̟ޟ���&�O� J�\�n���������߯ گ���'�"�4�F�o� j�|�������Ŀֿ�� ����G�B�T�fϏ� �ϜϮ���������� �,�>�g�b�t߆߯� �߼���������?�:�L�^����`l_INFO 1�i�` �U`��������
�?��@B?�z=��%�������A�m7�?	�_���?µ�B���k`YSDEBUGx`��`��d�i��SP�_PASSxeB�?��LOG v�e�a  ��9M���  ��a��UD1:\��<����_MPC���eHI[�ay �a~)SAV ��`�a������SV}�TEM_T�IME 1����` 0  �����{{���SKMEM  ��e�a�� %�{`rX|�`�(��� @��"����`�P�� ���b/ �`)�� �@�>/P/b/t/��/�B ��/����/�/�/�/��?? 1?C?U?g?y?�?�?�?Ike�?�?�?OO*O <ONO`OrO�O�O�O�O �O�O�O__&_8_�a�T1SVGUNS��`ye'�e�MPA�SK_OPTIO�Nx`�e�a�amQ_�DI��o�UBC2?_GRP 2;�c0��_6"0C��SA\�BCCFG ��[�(�!k8m`8o,�po[o�o�o�o �o�o�o�o�o6! 3lW�{��� ����2��V�A� z�e�������ʏ�� ������E�0�i�T� �����T����۟ɟ ���#��G�5�W�Y� k�����ů���ׯ� ���C�1�g�U���y� ��������ӿ	��ڀ �/�M�_�q�ￕσ� ���Ϲ�������7� %�[�I��mߏߑߣ� ��������!��E�3� U�{�i�������� �������A�/�e�� }���������O����� +OasA� ������� 9']K�o�� �����#//G/ 5/W/Y/k/�/�/�/{� �/�/??1?�/U?C? e?�?y?�?�?�?�?�? �?O	O?O-OOOQOcO �O�O�O�O�O�O_�O _;_)___M_�_q_�_ �_�_�_�_o�_%o�/ =oOomoo�oo�o�o �o�o�o!3W E{i����� ����A�/�e�S� u����������я� ����+�a�O���;o ����͟ߟ�o��� %�K�9�o�����a��� ��ۯɯ�����#� Y�G�}�k�����ſ�� տ�����C�1�g� U�w�yϋ��ϯ��ϛ� ���-�?�Q���u�c� �߫ߙ���������� �;�)�_�M�o�q�� ����������%�� 5�[�I��m������� ��������!E�� ]o���/�����/M�$�TBCSG_GR�P 2��  �M 
 ?�  x �t�����/��,/>+QX__d@ �m!?M	 HBL>(M�&~=$B$  C�p0�/�(}/�/Cz�/�-�A�>(333?&�ff?��<%A���/@?0 >(�1�a6&5V0DHC?�=@�0=%1�5=$�1D"!!�?�?[?�?O �:�(&�(AETOO1O O�OgOyO�O�O�K�H�Q	V3.0�0p	lr2d�C	*/P'TL>_f�O aQ�I uPG]v_  �_�_�[QJ2X_Q�_~�UCFG �i l�Z�rb�_Jn�Jo po~j"~o�o�o�o�o �o�o�o41j U�y����� ��0��T�?�x�c� ������ҏ������ ,�p� 7�I�[���� y���ğ���ӟ��� 0�B�T�f�!���u��� �����M9	�� �-�c�Q���u����� Ͽ��߿��)��M� ;�q�_ρσϕ��Ϲ� ������7�%�G�m� [ߑ�ߵ��߇���� ���3�!�W�E�{�i� �����������	� ��S�A�w������� g��������� O=sa���� ���9'] Kmo����� ��#//3/Y/�q/ �/�/?/�/�/�/�/�/ ??C?1?g?y?�?�? [?�?�?�?�?�?O-O ?O�?OOuOcO�O�O�O �O�O�O�O�O_;_)_ __M_�_q_�_�_�_�_ �_o�_%ooIo7oYo [omo�o�o�o�o�o�o �/'�o�oiW� {������� /��?�e�S���w��� ��я㏝����+�� ;�a�O���s�����͟ ��ݟߟ�'��K�9� o�]�������ɯ��� ۯ���5�#�E�G�Y� ��	����˿u���� �1��U�C�y�gϝ� �����ϑ������	� +�Q�c�u�/�A߫ߙ� �߽�������'�M� ;�q�_������� ������7�%�[�I� �m������������� ��!3ݿK]� ������� ASe#5�� ����//�=/ +/M/O/a/�/�/�/�/ �/�/?�/?9?'?]? K?�?o?�?�?�?�?�? �?�?#OOGO5OkOYO {O�O�O�O?q�O_ �O�O_1_g_U_�_y_ �_�_�_�_�_	o�_-o o=o?oQo�o�o�o�o wo�o�o�o)9 ;M�q���� ���%��I�7�m� [�����������ُ ���3�!�W�i�_�� ����O�՟ß���	� ��S�A�w��������k�ѯ������� s ?�C� C��W�C��$TBJO�P_GRP 2 ��� / ?�C�	o�v��"}�����@� �0��  � �� � � �=C� @?���	 �BL  �?Cр D]��������&�<��B$鰌��@���?�33C���X��f�q���x'ϩϷ�;�2�G�����@��?����z��_� �A��ȍ�� �Ϡ����?�>�Q�4�F�;���pA��?�ff�@&ff?�ffWψ�� ��ߝ�P�x������:v,���c?LQ�P�t�DH��x�� �@�333儯���>t�O�X�j�8����3Ꮁ���D"�������3�E�O�x������9���� ��:�I�T�K���s�]� k�������_����� ��)Z5��y�}0���C�C�C�ܱ���	V3.0~Ƴ	lr2d���*5��>�CN� E8� EJ�� E\� En�@ E��E�� �E�� E�� �E�� E�h �E�H E�0 �E� E�e��� E�i� �E�x E�X �F�^D�  �D�` E}�P Ee$m0��;iGqR�^op Ekyu�rڥ���(z� �E�}���X O9�IR!�%�
M�3/E"C��I#��߄/k�ESTPARS 7���l��HR� ABLE �1#}� C�D�(^' ��>)�'�(��(B�J��'	�(
��(�(�%C��(�(�(!�#RDI�/���/�/�/??15�4O�?�;�?�?�?H�?N�"S�?�� c: �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oob��@�O�� �']iFOXOjO|O(?:?�L?^?p?�8�"CbNUoM  ���ϰK�   �"_CFG $,{��c�@o�IMEBF_TT�!�e��� �nvVER#oa�v�nsR 1%�+ �8@C�>��q �ho  ���� �#�5�G�Y�k�}��� ����ŏ׏����V� 1�C���g�y������� ��ӟ���	��-�?� Q�c�u���������ϯ ���N�)�;���_� q���������˿ݿ�"R�q_&q�v@�u� MI_CHANzw� �u H�DBGL�V��|u�u�!K�E�THERAD ?U�%���I ��￷��ϓ(K�ROUmT�p!*J!������SNMASK��ȥs��255.�Y�!W�i�{�!� O�OLOFS_DI� �}�ORQC?TRL &�{CJ/��T���/�A�S� e�w��������� ����+�=�M���p��_����#PE_DE�TAIqȾ�PGL�_CONFIG �,,y<q��/�cell/$CID$/grp1��@ 2DVC��� ������j� #5GY�}� ����fx// 1/C/U/g/��/�/�/ �/�/�/t/	??-??? Q?c?�/?�?�?�?�?�?�?gn}�?)O;OMO�_OqO�O�a���O�M� �?�O�O__(_:_�? ^_p_�_�_�_�_G_�_ �_ oo$o6oHo�_lo ~o�o�o�o�oUo�o�o  2D�ohz� ����c�
�� .�@�R��v������� ��Џ_����*�<� N�`��������̟ ޟm���&�8�J�\� 럀�������ȯگ����User� View ��}�}1234567890�/�A�S�e�`w��������2�|�����)�;Ϛ���
�3Ŀ�ϛπ�Ͽ�����B�߲�4 x�=�O�a�s߅ߗ����߲�5,�����'� 9�K��lﲾ6�ߥ� ����������^� ���7��Y�k�}������������8H�1�CUg���� �lCamera����'BE�Qcu ���������  �ù�9/K/]/ o/�/�/:�/�/�/&/��/?#?5?G?Y?�� �w��/�?�?�?�?�? �?�/#O5OGO�?kO}O �O�O�O�Ol?~7+�\O _#_5_G_Y_k_O�_ �_�_�O�_�_�_oo 1o�O~7+�_o�o�o �o�o�o�_�o!lo EWi{��Fo� ��4����1�C� �og�y��������ӏ ���	��~7G���U� g�y�������V�ӟ� ��B��-�?�Q�c�u� �~7�����ӯ��� 	��?�Q�c������������ϿῈ���9 m�"�4�F�X�j�|�#� �ϲ���k�������P0�B�T���	�0�� �ߡ߳������ߐ�� �1���U�g�y��� ��V�h߮ �S��� ,�>�P�b�	������ ��������(�� �+��t���� �u��a:L ^p��;uՈ;+ ��//(/:/�^/ p/�/��/�/�/�/�/  ?���K�/L?^?p? �?�?�?M/�?�?�?9? O$O6OHOZOlO?� `kO�O�O�O�O __ �?6_H_Z_�O~_�_�_ �_�_�_O��{o_$o 6oHoZolo~o%_�o�o �oo�o�o 2D�]  �Ys� ��������<'�9�   IQ o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u�������=��  
�P(  }�gp( 	 �� �߿��9�'�]�K� m�oρϷϥ�������:źY� ̓oD� V�h��o�ߞ߰����� ���S3��"�4�{�X� j�|���������� ��A��0�B�T�f�x� ������������ ,>����t�� ������] :L^����� ��# //$/kH/ Z/l/~/�/�/���/ �/�/C/ ?2?D?V?h? z?�/�?�?�?	?�?�? 
OO.O@O�?dOvO�O �?�O�O�O�O�O_MO _O<_N_`_�O�_�_�_ �_�_�_%_oo&om_ Jo\ono�o�o�o�_�o �o�o3o"4FX j�o�o���� ���0�B��f�x� �������ҏ���� O�,�>�P���t�����ટ��Ο���@  ����!����۰���+frh:\�tpgl\rob�ots\lrm2�00id[�_ma�te__�.xml ݟ��������ϯ��0��)����3�X� j�|�������Ŀֿ� ����5�/�T�f�x� �ϜϮ���������� �1�+�P�b�t߆ߘ� �߼���������-� '�L�^�p����� ������ ��)�#�H� Z�l�~����������� ����%�DVh z������� 
!@Rdv� ������/.::�p� ��E��<< C� ?�+[//S/u/�/�/ �/�/�/�/?�/?)? W?=?_?�?s?�?�?�?�?�?O��$TP�GL_OUTPU�T /#�#� ; CEXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_CE; ��@2345678901o-o?oQo couo}c�o�o�o�o �o�o�o�o4FXj|z}���� ����,�>�P�b� t��������Ώ��� ����:�L�^�p��� �,���ʟܟ� �� �� �H�Z�l�~���(� ��Ưد�������� D�V�h�z�����6��� Կ���
�ϴ�*�R� d�vψϚ�2�D����� ����*���8�`�r� �ߖߨ�@߶�������&��A}6!\�n� �������@=/�����C* ( 	  o2� �V�D�z�h� �������������� 
@.dRt�� ����� *`N�f�9 R& �����/�(/ :/j�k/}//�/�/ �/�/�/�/Y/�/1?�/ ?g?y?S?�?�??�? �??�?O-OOQOcO �?KO�O�OEO�O�O�O �O_uO�OM___�Og_ �_o_�_�_�_;_oo �_�_Io#o5oo�o�_ �o�oao�o�o�o3 E�o-{�'�� ���W�/�A�� e�w�Q�c������ �����+���a�s� яw���C���ߟ�˟ �'����]���I��� ���ɯۯ9�ï�#� ��G�Y�3�e������ ſ׿q�߿����C� Uϳ�yϋ�%�w��ϛ�����	ߛ�$TP�OFF_LIM ���М����$�N_SV(� � ��:�P_M�ON 0��<�����2��$�S�TRTCHK �1�:�Y�B�VT?COMPATO����>�VWVAR �2o���S� R�� �3���$��_DEFPROG� %��%-BCKEDT-+����_DISPLA�Y/О�D�INST�_MSK  ��� ��INUSE9R�߆�LCK����QUICKMEN����SCRE�����tps�c����6�;�:�L�_�P�ST��:�RAC�E_CFG 3�o���3�	�
�?���HNL 2!4S�x��� )��� %7I[m
���ITEM 25��� �%$12�34567890<��  =<��<  !&��_���� ���>P/t 4/�D/j/���/ /(/�/L/�/?0?�/ T?�/�/�/V? ?�?�? �?H?�?l?~?�?ObO �?�O�O�?�O O2O�O VO_zO:_L_�Ob_�O &_�_
_�_._�_ oo v_o�_�_�_8o�_�o �o�o*o�oNo`oro�o �ohz�o� �8�\�.��D� ����������� h�X�j�|������ď p������̟0�B�T� Οx�$�J�\���h�� �����گ>����t� �����s�ί��򯲿 Ŀ(�ڿL���'ς�B� ��R�xϊ���$� 6ϰ�Z��,�>ߢ�b� ������n߆� ����� V���zߌ�U��p��� ���
��.�@�	����S��6���� 3 �� ��e�\�
 r������~=�UD1:\����� �R_GRP� 17�� 	 @e�&@F4jX�|��  ��
������?�  ,>(^ L�p�����  /�$//H/6/l/Z/|/�/	��/�/�SCB 28*� ?&?8?J?\?�n?�?�?�?�UTORIAL 9*�����?�V_CON?FIG :*����b���NO�=OUTP�UT ;*�?@��ZO�O�O�O�O �O�O
__._@_R_d_ v_<A�O�_�_�_�_�_ �_
oo.o@oRodovo �_�o�o�o�o�o�o *<N`r�o� �������&� 8�J�\�n�������� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t��� ������ο���� (�:�L�^�pςϓ��� �������� ��$�6� H�Z�l�~ߏϢߴ��� ������� �2�D�V� h�z��(O:E�O���� �� ��$�6�H�Z�l� ~���������������  2DVhz� �������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/��/ �/�/??&?8?J?\? n?�?�?�?�/�?�?�? �?O"O4OFOXOjO|O �O�O�O�?�O�O�O_ _0_B_T_f_x_�_�_ �_�O�_�_�_oo,o >oPoboto�o�o�o�_ �o�o�o(:L ^p�����o� � ��$�6�H�Z�l��~������������ӏ�ρ����� 4�F�X�j�|������� ğ֟�����0�B� T�f�x���������ү �����+�>�P�b� t���������ο�� ��'�:�L�^�pς� �Ϧϸ������� �� #�6�H�Z�l�~ߐߢ� ����������� �1� D�V�h�z������ ������
��-�@�R� d�v������������� ��)�<N`r ������� &7J\n�� ������/"/ 3F/X/j/|/�/�/�/��/�/�/�/??-;��$TX_SCRE�EN 1<��π�}i�pnl/a0gen.htm-?�?�?�?��?�?%�Pan�el setup�<}��?OO1OCOUOgO�?�?�O�O�O �O�O�OoO_�O@_R_ d_v_�_�__#_�_�_ �_oo*o�_�_�_ro �o�o�o�o�oCo�ogo &8J\n�o�o ������u� �F�X�j�|������ ď;������0�B����0>UALRM_�MSG ?M9�Z0 [�0*����؟ ˟��� ��%�C�I��z�m�����¯v�SEoV  �����t�ECFG >vM5W1  0%�@�  A$�  w B�0$
 ï 7#M5W�i�{��������ÿտ����� �G�RP 2?
� 00&	 A�c�v��I_BBL_NO�TE @
�T?��l7"R0�9!�v�DEFP�RO��%�� (%����9 �����(� �L�7�p�[߁ߦߑ���ߵ���l�FKEYDATA 1AM9�M�p �0& �R�d��A����w�,(����0$��|����ANCEL��-���Q�8�EXT STEPZ�]��������ORE INFO��������( L^E�i������  ���  frh/gu�i/whitehome.png Qcu��(������//�FR�H/FCGTP/�wzcancel <V/h/z/�/�/��/��/�/�/
??'/9#nextE/\?n?�?�? �?�/�?�?�?�?O"O<-?7#infoK?bO tO�O�O�O�?�O�O�O __(_�OL_^_p_�_ �_�_�_G_�_�_ oo $o6o�_Zolo~o�o�o �oCo�o�o�o 2 D�ohz���� Q��
��.�@� O�v���������Џ� ���*�<�N�ݏr� ��������̟[�ޟ� �&�8�J�\�럀��� ����ȯگi����"� 4�F�X��j������� Ŀֿ�w���0�B� T�f����ϜϮ����� ��s����,�>�P�b� t�ߘߪ߼������� ���(�:�L�^�p��� ���������� ���$�6�H�Z�l�~�U�����$���������������,�=�aH�� ~������ 9K2oV��� ����/#/
/G/ ./k/}/\��/�/�/�/ �/�/
�?1?C?U?g? y?�??�?�?�?�?�? 	O�?-O?OQOcOuO�O O�O�O�O�O�O__ �O;_M___q_�_�_$_ �_�_�_�_oo�_7o Io[omoo�o�o2o�o �o�o�o!�oEW i{��.��� ���/��S�e�w� ������<�я���� �+���O�a�s����� �����/ߟ���'� 9�@�]�o��������� ɯX�����#�5�G� ֯k�}�������ſT� �����1�C�U�� yϋϝϯ�����b��� 	��-�?�Q���u߇� �߽߫�����p��� )�;�M�_��߃��� ������l���%�7� I�[�m���������� ����z�!3EW i����������А��А���$6H j|V,h/�`/� ��/�+//O/a/ H/�/l/�/�/�/�/�/ ??�/9? ?]?D?�? �?z?�?�?�?�?̟O #O5OGOYOkOz�O�O �O�O�O�O�O�O_1_ C_U_g_y__�_�_�_ �_�_�_�_o-o?oQo couo�oo�o�o�o�o �o�o);M_q ������� ��7�I�[�m����  ���Ǐُ������ 3�E�W�i�{�����.� ß՟�������A� S�e�w�����*���ѯ �����+�OO�a� s���������Ϳ߿� ��'�9�ȿ]�oρ� �ϥϷ�F�������� #�5���Y�k�}ߏߡ� ����T�������1� C���g�y������ P�����	��-�?�Q� ��u�����������^� ��);M��q ������l %7I[�� ����h�/!/�3/E/W/i/@�k+}�@�����/@�/�-�/�/�/�&,�? ?�?A?(?e?w?^?�? �?�?�?�?�?�?O+O OOO6OsO�OlO�O�O �O�O�O_�O'__K_ ]_<��_�_�_�_�_�_ ��_o#o5oGoYoko �_�o�o�o�o�o�oxo 1CUg�o� �������� -�?�Q�c�u������ ��Ϗ�󏂏�)�;� M�_�q��������˟ ݟ����%�7�I�[� m�������ǯٯ� �����3�E�W�i�{� �����ÿտ���� ��/�A�S�e�wωϛ� r_���������� � =�O�a�s߅ߗߩ�8� ��������'��K� ]�o����4����� �����#�5���Y�k� }�������B������� 1��Ugy� ���P��	 -?�cu��� �L��//)/;/ M/�q/�/�/�/�/�/ Z/�/??%?7?I?�/ m??�?�?�?�?�?����;������OO(M OJO\O6F,H_�O@_�O�O�O �O�O_�O/_A_(_e_ L_�_�_�_�_�_�_�_ �_o o=o$oaosoZo �o~o�o�o���o '9KZ?o��� ���j��#�5� G�Y��}�������ŏ ׏f�����1�C�U� g�����������ӟ� t�	��-�?�Q�c�� ��������ϯ�󯂯 �)�;�M�_�q� ��� ����˿ݿ�~��%� 7�I�[�m��ϣϵ� �������ό�!�3�E� W�i�{�
ߟ߱����� ������o/�A�S�e� w��߭�������� ����=�O�a�s��� ��&��������� ��9K]o��� 4����#� GYk}��0� ���//1/�U/ g/y/�/�/�/>/�/�/ �/	??-?�/Q?c?u? �?�?�?�?L?�?�?O O)O;O�?_OqO�O�O �O�OHO�O�O__%_h7_I_ �K[� ����t_�_�]p_�_�_�V,�o�_�o !ooEoWo>o{obo�o �o�o�o�o�o�o/ SeL�p�� �����+�=�� a�s����������Oߏ ���'�9�K�ڏo� ��������ɟX���� �#�5�G�֟k�}��� ����ůׯf����� 1�C�U��y������� ��ӿb���	��-�?� Q�c��ϙϫϽ��� ��p���)�;�M�_� �σߕߧ߹������� ~��%�7�I�[�m��� ����������z�� !�3�E�W�i�{�R��� ���������� �/ ASew��� ����+=O as����� �//�9/K/]/o/ �/�/"/�/�/�/�/�/ ?�/5?G?Y?k?}?�? �?0?�?�?�?�?OO �?COUOgOyO�O�O,O �O�O�O�O	__-_�O Q_c_u_�_�_�_:_�_ �_�_oo)o�_Mo_o@qo�o�o�o�o���k���������o�o}�o*<v, (�m ��x��� ���!��E�,�i� {�b�����ÏՏ���� ����A�S�:�w�^� ������џ����� +�:oO�a�s������� ��J�߯���'�9� ȯ]�o���������F� ۿ����#�5�G�ֿ k�}Ϗϡϳ���T��� ����1�C���g�y� �ߝ߯�����b���	� �-�?�Q���u��� �����^�����)� ;�M�_���������� ����l�%7I [������� �!3EWi p������� �///A/S/e/w// �/�/�/�/�/�/�/? +?=?O?a?s?�??�? �?�?�?�?O�?'O9O KO]OoO�OO�O�O�O �O�O�O_�O5_G_Y_ k_}_�__�_�_�_�_ �_o�_1oCoUogoyo �o�o,o�o�o�o�o	 �o?Qcu�� (������)�� +�� ���T�f�x�P�������,��ݏ���� %�7��[�B����x� ����ٟ�ҟ���3� E�,�i�P���t���ï ���ί���A�S� e�w��������ѿ� ����+Ϻ�O�a�s� �ϗϩ�8�������� �'߶�K�]�o߁ߓ� �߷�F��������#� 5���Y�k�}���� B���������1�C� ��g�y���������P� ����	-?��c u�����^� );M�q� ����Z�// %/7/I/[/2�/�/�/ �/�/�/��/?!?3? E?W?i?�/�?�?�?�? �?�?v?OO/OAOSO eO�?�O�O�O�O�O�O �O�O_+_=_O_a_s_ _�_�_�_�_�_�_�_ o'o9oKo]ooo�oo �o�o�o�o�o�o�o# 5GYk}�� ������1�C� U�g�y��������ӏ ���	���-�?�Q�c��u�����p ���>p ���ğ֟ ���
����,�M�  �q�X�������˯�� ���%��I�[�B� �f�������ٿ���� �!�3��W�>�{ύ� l/������������ /�A�S�e�w߉ߛ�*� �����������=� O�a�s���&���� ������'���K�]� o�������4������� ��#��GYk} ���B��� 1�Ugy�� �>���	//-/ ?/�c/u/�/�/�/�/ L/�/�/??)?;?�/ _?q?�?�?�?�?�?�� �?OO%O7OIOP?mO O�O�O�O�O�OhO�O _!_3_E_W_�O{_�_ �_�_�_�_d_�_oo /oAoSoeo�_�o�o�o �o�o�oro+= Oa�o����� ����'�9�K�]� o��������ɏۏ� |��#�5�G�Y�k�}� �����şן����� �1�C�U�g�y���������ӯ���	��$�UI_INUSE�R  ����*�� � 
��_MENHIST 1B*��  �( 7���(/�SOFTPART�/GENLINK�?current�=menupage,153,1I�p��ο��� ����962��>�P�b�0t���'�36-��� �����χϙϫ�@�R� d�v�ؓߥ߷����� ���ߎ�#�5�G�Y�k� }������������ ���1�C�U�g�y�������~�������� ���9K]o ��"����� ��GYk}� �0����// �C/U/g/y/�/�/,/ >/�/�/�/	??-?�/ Q?c?u?�?�?�?���� �?�?OO)O;O>?_O qO�O�O�O�OHO�O�O __%_7_I_�Om__ �_�_�_�_V_�_�_o !o3oEo�_io{o�o�o �o�o�odo�o/ AS�ow���� ��?�?��+�=�O� a�d��������͏ߏ n���'�9�K�]�o� ��������ɟ۟�|� �#�5�G�Y�k����� ����ůׯ������ 1�C�U�g�y������ ��ӿ�����-�?� Q�c�uχϊ��Ͻ��� ����ߔϦ�;�M�_� q߃ߕ�$߹������� ���7�I�[�m�� �� �2���������� !���E�W�i�{����� .�������������$UI_PA�NEDATA 1�D���S�  	�}�  FRH/FC�GTP/FLEX�UIF.HTM?�connid=0�/�����) � rim��   d $6HZl� ~�������  //D/V/=/z/a/�/p�/�/�/�� ��"	? ?2?D?V? h?�/�?��?�?�?�? �?
OO�?@O'OdOKO vO�O�O�O�O�O�O�O�_�O<_N_5_r_�, �VU�?�_�_�_�_�_ ob_3o�?Woio{o�o �o�oo�o�o�o�o /A(eL�p� �������_�_ O�a�s��������͏ @o���'�9�K�]� ď��h�����ɟ۟ ���#�5��Y�@�}� ��v���&�8����� �1�C���g�y�쏝� ����ӿ���^��� ?�Q�8�u�\ϙϫϒ� �϶������)��M� ��ү���ߧ߹����� ��B�7�I�[�m� ���ߵ�������� �!��E�,�i�P��� ������������l�~� /ASew����  ����+= �aH�l��� ��//�9/ /]/ o/V/�/�/�/�/ �/?#?v/G?Y?�}? �?�?�?�?�?>?�?�? O1OOUO<OyO�OrO �O�O�O�O�O	_�O-_�/�/}�>_w_�_�_�_�_�_)e_�_i5�_ "o4oFoXojo|o�_�o �o�o�o�o�o�o BT;x_�����b8�#�+�$UI�_POSTYPE�  �%� 	 �5���QUICKMEN  �"�8���RESTORE �1E�% � ��k2������k2mڏ�� '�9�K��o������� ��Z�۟����#�Ώ 0�B�T�Ɵ������ů ׯz�����1�C�U� ��y���������l�ο ��d�-�?�Q�c�u� ϙϫϽ����τ�� �)�;�M����l�~� �Ϣ���������� 7�I�[�m��"��� ���������
���� W�i�{�����B����� ������ASexw�C�SCRES��?X�u1�sc��u2�3��4�5�6�7r�8��TAT��� g��%�zUS#ER� ��T� �Sks�_4_5_�6_7_8_�N�DO_CFG �F�NPMQ�OP_CRM5  IU���PDA�NoneF��8_INFO 1�G�%	 e�0% �$/b8/S/6/w/�/ l/�/�/�/�/�/??��/=?O?2?s?<��O�FFSET J�!�?*��2�? �?�?�?'OO0O]OTO fO�?jO�O�O�O�O�O �O#__,_>_�Kh��]�x_�_
�_�_�8UF�RAME��SR�TOL_ABRT8�_�bENBoh?GRP 1K��d�Cz  A�mc ka,ko}o�o�o�o�f!�o�ojR�U7h�~&kMSK  :e�	!&kN�Q%)��%Z_{E�VARS�_CONFI�Ln�; FP*��x�CMRSb2R�;y, 	��p`0�1: SC13?0EF2 *�
�J*�OX��t��[ �?��`@�`up�`�~ �_^�h�#����ȏ�qhÏ��a��eA�,�܏-�, B���H�,L�ԏm� ����`�����ٟğ�� ���3����i�T�f����R�ïկ�tISI?ONTMOU`:t���쥙S�S��S�0�ba FR:\��\�A\گ �� UD1-�wLOG:�  S��EX_�,' ?B@ ����r��j��r�ÿ�* �� n6  ����#��t��`����  =����5�*2�s�TR�AIN����D¿P  dy�p5�"��
�rT�=(��5Ž�V� ����������4�"�8� F�X�j�|ߎߠ���W�Z�_��RE�UZi��r�tLEXE�V̡|�1-��~MP�HAS	���D��sRTD_FILTER 2W�; �RU�U���� ��������&�8�J� �J��{�����������������vSHI�FTr1X�;
 <��iwV| ������!� 
0i@R�v����	LIVE�/SNA�s%v�sfliv;���+� �0U�p
"menu /%/��/�/m"6�YE	Gr2�MO�Z'���`��$WAITDINGEND��#x�$O7p�7��*?S>?9T�IM8u��i<G �/�=?�;=?�:\?�:<{?8RELER�8o��$����!_ACT��=HCxrB6� [�\{�/�O�VrBRDI�S�p9o�$XVR��\'��$ZA�BCSc]� ,r�X2�O�]ZIP�^����_�_�_�TZMPCF_G ;1_Zk 0s�~_�o�WSc`Zi@q�� �茯Ro�a< +�Wo�o�oAo�oeiH� ���o�o�o�o�oA�ot�D��I��������{P�P�a�j_SbPYLIND�x�b�[ � �,(  *\�m���Y�0��}����� o�� ��V�7���[�B�T� ��ԏ��ǟٟ����� ~�3��W�>��������S[ c2c�W�A ��_����n#���G�Kyگw�Kw���A��*�SPHERE 2d<���ͿA� ƿ��'�o���]�o� 럓�2���ϰ����� F�#�5�|ώ�k��Ϗ� v߈���������PZZ\F �HF