��  	w^�A��*SYST�EM*��V9.1�0185 12�/11/2019� A  �����AAVM_�WRK_T  �� $EXP�OSURE  �$CAMCLB�DAT@ $PS_TRGVT��$X aH]ZgDISfWg�PgRgLENS_CENT_X��YgyORf  � $CMP_G�C_�UTNUM�APRE_MASwT_C� 	��GRV_M{$�NEW��	ST�AT_RUNAR�ES_ER�VTSCP6� aTCb32:dXSM�p&&�#END!�ORGBK!SMp��3!UPD�O�ABS; � P/ �  $P�ARA�  ����AIO_wCNV� l� �RAC�LO�M�OD_TYP@F+IR�HAL�>#�IN_OU�FA�C� gINTER�CEPfBI�I�Z@!LRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� �!PCOU�PLE,   �$�!PPV1CESI0�!H1�!"PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W� @V�R!SBN_�CF�!�0$�!J� ; 
2�1_C�MNT�$FL�AGS]�CHE�"$Nb_OPT��2 � ELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1 UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t�cbMO� �sE 	� [M�s��2�wREV�BILF��!XI� %�R 7 � OD}`j��$NO`MD�+� `�x�/�"�u�� ����^��@D�d p E R�D_Eb��$F�SSB�&W`KBD�_SE2uAG� G
�2 "_��B�� V�t:5`ׁQC���a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR��BIGALLOW� (KD2�2�@VAR5�d!�A>B ��BL[@S � ,KJqM�H`9S�pZ@M_O]z�ޗ�CFd �X�0GR@��M�NFLI���;@UIRE�84�"� �SWIT=$/0_N�o`S�"CF_�G�� �0WAR�NMxp�d�%`LI��V`NST� CO�R-rFLTR^�TRAT T�`>� $ACCqS��� X�r$ORIأ.&ӧRT�`_SYFg��HGV0I�Ep�T��PA�I��5T���HK�� � �#@a��N�HDR�B��2�B�J; �C��3�4��5�6�7�8�  �0��x@�2� @� TRQB��$%f��ր����c_U���� COc <� ����Ȩx3�2��LLECM�}-�MULTIV4��"$��A
2FS�I�LDD��c� DET}_1b  4� STY2�b4�=@��)24��e`DԼ� |9$��.p��6�aI`�* \�TO�:�E��EXT����p���B�ў22�0,D��@��1b�.'�B ��G�Q� �"Q�/%�a��X� %�?sdaD�U� Sҟ؈;A�Ɨ�M�� �� CՋO�! L@�0a�� X׻pAβ$JOBB���֍�v��IGO�" dӀ �����X�-'x���G��ҧ]�C�`��b# etӀF� �CNG�AiBA� ϑ��!��� /1��À�0����R0aP/p3���$
��|��BqF]�
2J�]�_RN��C`J�`�e�J?�D/5C��	�ӧ��@����Pr�O3л!% \�0�RO�6� �IT<�s� NOM_8pn#��c ���TU��@P� � ��&"+P��� ӨP�	ݭ��RAx@n �3�A����
$TF3%#D%3
T��wpU�13��}�%mHrzT1�E���ޣ�#ݤp�%ߢQlYNT�"�� DBGDE�!'D�]�PU���@t����"��AX��"�uwTAI2sBUFۆ;%�1( ��P&V`[PI84'mP�'EM�(M�)B �&F�'�SIMQS�@ZK;EE3PAT�z�`�8"�"�MC��1)S�0��`JB�����aDECg:� g5e������* �U�CH�NS_EMPͲ#$G��7�_��c�;�1_FP)�TC�6S���5�`%��4�} ��V����W���JR����SEGF�RAq�O�� #PT�_LIN�KCPVAF���`  C$+�� �ckBZ��PBzr���@>6,` +�Ԧ ��A�0��Ad0o`Arp�D���Id1SIZh���	T�FT�C�Z1Y�ARSm��CP@'�@Ic\1@cX�0<@L��8��0�VCRCߥ�sCC���U1@�X�1��2�Mpq�U�1`�XD�Q�UDݤأiCk �p��
DK`݀f��RhSEVRf �Fha_	EF�0N�f�Pd1�&hB��5�jC}�+�OVSCA[��A�f����13��-�	<�ׇMARG���"a�F@@���1DcQ�rN�0LEW�-��R��P<��o�l��RɄ.� ����ǯ��� 5ڡR�`HANC��$LG5��a��Ӑ��ـF��Ae����0RYr�3
����
��@ �RA��
�AZ��0Q�N`�O��FCT��sp�F��R�0\P0b ADI��O�� +���+���&���5�5Є���S[�g���BMPUD(PY�1��GAESCPjc��W��%N  S-��U0ۑuU�/)�TIT'q�<�b�%ECA:!�!E'RRLd��0�&Q��OR�B$������~Ұ$RUN_O��SYS��4������u�REV�V@��?DBPXWO�P�=10�$SKo�"�1�DBT�pTRLn�2 �C AC��0��%�m�U DJ�p��_�`�!A�ǀM�P5L�A_2WA��j�EE��D!w�!%R|hO�UMMY9��ڠ�1� ��DBd[��3���!PR�Q� 
��ٱ9��4� г$r��$ Q��Lة5L�z����6�^z�PC�7*��<�ENEC0Tq�8I�����RECO}R$�9H mގ�4$L��5$ أ�"E���R@��VA��s_Dց� ROS �"SK�����I�=�א��PA��JVB�ETURN���SMeR(�U #�CRʰ�EWMDB0GNsALV �"$LA� �[�*6$P-�g7$Pv�s�8o��!�PC��#�DO�^@-�Ŵ���R˶GOg_AW�ܱMOz���p���CSS_+CN4�YO�:��T���0���ID�T�2*��2�N��O@�J���v`Iְ ; oP $>�RB�B���PI�POl�IG_BY��vЅ�TVR���HNDG$�< H�`�1a�@cS��DSBLI��s��ְ0}����LS$�=0��0� ��FB�FEձL�9����5z��>D�$DO�1�C�pMC�0q��4(��9�RH��W��K�4ELE�ur�
^��SLAVr?xB�INS ���#����_R@P�@\`�pS� }�l�}�l�{u��[!e��ے�I���B�r�W��D�NTV�#��VE�$��SKI lA4;3��2UB�1�J�f�1C�
DSAF�7�5��_SV6�EOXCLU-��Xr'ONL�0YY��s<����HI_VՀ�R�PPLYo�RCsHX� �0_M�QПVRFY_I�.Mms$IOv0��}"��1UB���Oj�3�LS����4!���:@�P�$��ĆAUTOCN�E ����.��GCHD�s��_���3sЛAF��CPe�T�!��р� A�o���_�0  �Ԣz�NOCtB$xB�pT��A �����SG�` C� � 
$CUR 8�U��!" �� T@B������ANNUNC�#���䱐b���()%!��-*I&��p@��IC�D @b�`F
"a��POTX� aө�����������[EM��NIߢE��ȷ"�G� A��$DA=Y��LOAD`Ԟ���"��5�� �EF_F_AXI�Fo��%Q�O0<�:�_�RTRQV1G D�a��?0�RK3�0S45 2Fz@]w:1�a�d�A0p/1sAH 0B!�1A�T�2�æ�vDUX��u��C�ABsAIs"�pNSl�1�PID�@PWSsh�5�AWpV`�V_�0|q0�P�DIAGy�sAJ� 1$VX��ET	`�UrT��EJā�{RRf��!�TVE6�� SW|AZ� sP�0�:5q0G}P:13OHP5�1PP|@�SIR|�{RB�P�2�3 %qZQC �BB��H� ^��E`��5q0I��?0����URQDW�EM	SB�?UA�p�EjB�TLIFE�`K#iP��uRN|QFB�U%!zSFBh�a�%"C����N��Y'p�FLA��t& OVڰ�VHE|��BSUPPO(��uRI�_�T��QC_X�d�� gZjWj� g��%!��6�cXZ*�ϡfAY2xhEC��T��DEN�pTBE%!J�� �F_8p��A� @CT�K{ `Q�CACH�*r�bSIZ�V�Pz`�N��UFFI`�oP�ឤ2���62��M;��tL �81 KEYIMAG �TM��!�^q:��Yv�����OCVI9E�@�qM �༠�L~��;�?� 	���р�dNG0��ST��!�r���t����t0�t0�pEMA�ILo����!�5FAUL�"O�r��/����COU��쑁�T���)AP< $d9�p�S�0�0IT��BUF�g;��gE�o�Je��PBe�p�C:�p��:�|�G�SAV�� r�[@�b��@ˇÐ)&AP��p印�D��_e���� �OT겮�3�Pm ��0�z3�AX��#f x Xe�C�_uG|S
^YN_�A.��Q <I0Dk�O�����BM�2�PT�� F!�$�D�I[E7�����R$��$ G���!&�Ǳད�:�9�S�0���-��C_ᰤ�AK�$�����RVq8���DSPnv�PCe�IM��\���<�3@U9��P�] �IP���A�`[�CTH�`3�O�0T��\�HSȓ>�BSC���`e�V��
��#X���*4NV��G;����`Y�e�F|A}�d0>���Z�"�SC%Ba���MER)�FBgCMP)�ET�� TLrFU`D�UY���R�mb�CD R�ܠ'�"���R��
n!UG0*����%��R�%P���C�
ń�-"2��:�o V/H *
�L�� )�9���G ���}�Z {ƥ!{�1{�1{�6q*{�7x�8x�9x�|PTzȄ�1��1��1��U1��1��1��1�ʕ1��2��2�ˑ�2���2��2��2��2���2��2��3��3R��3�˞�3��3��U3��3��3��3��94��61EXT6An!W��߸���V��uş�t���@FDR%D/XTE�V� .�puR�
�uRREM^@9F���BOVM5�*��A3�TROV3�D�T��S�MXb�INp3��PR�"AINDq�BcB
��ɐ}���Ge� �C\�p�UkADO6\��RIVW�R�BGE[AR5�IObEK#�cDN��1`X� zp|`dCZ_MCMp`nuQ �F�PUR���Y ,���?� �P>?o {A?oE� w�1�������Z0*PPM��2@RI��r�ET�UP2_ [ �0q�TDʠ�1p�T�����5�r�BAC��\ T�pr�蔅)�%w#@ó�TIFI�A����d��@/�PT�B�FLUI�t] �@�x;�UR�A���R�Б
���:C_0I�$�S�_?x�J�C9O��"�VRT��� x$SHO^14 #�ASS�-��U̠��BG_ �!.�!���!��!��FORCz#��hDATA)A-^�rFUZ1��]#�2��ˑi�`)A_ �|��NAV=�)�����S��S?$VISI��SC=�SE� ��5UV� O�1&1BFx�4@�&$PO� �I�A�FMR}2��` � ��2���6�!�3J�)�CE#�_����_@IT_Yִ]@�M������DGCL�F�EDGDY�8L�D���5�V���TRH M���sa4�v9? T�FS
��t�b P��RB��}��$EX_RAiHRA1PY�X��RS@3�K5�Fs�G&�	5c �� ֳ�SW��O0VDE�BUG$�A(�GRt� opUz�BKU���O1M� �0P�OZ0Y�@���E�@M��LOOM�9QSMz�0E�� d�����P_E d x�P���TERM[UyedU��ORI֑�`PfdUa0�SM_��`Pg�V�`Q �X�hdU��UP�rig� -���2d��rS�Pe� G�Z @E�LTO���A�FIG�bZ �Agp�T��Tf$UFR��$��aM`ѵ�0OTZgA�TA��lcwNSTאPAT�<�`�bPTHJ�ϰ�E�p�ذbART�؀"e)�؁���REyL�j�SHFTӢ(�a�h_�R��̳J�V �P$�Wph�1p����t�SHI�`�4U � ҁAYLO��m���l� ��a8}!�ޠERV��Sq �x��hgא�b �K��u.�KRC��A�SYM���WJ+g���E��a�y�ұU�א���e@�v��eP��ppE�2vOR2אM3� GRJQ
4jX"�B0V�`G`l�� sHO�6Dk ��aXN� �OCaQ>@$OP�$e��i�����d�ՀRY��aOU��c�PTR�e���|�a�e$PWR��3IM��rR_˃�d0� �P�cUD��c�SV򳠁֔l� �$H�!��ADDR��HMQG�b����ʨ���R�"1m H��S���! ��.�0畞�畫�SEz1�#�PHSܰ
3n $Z À_D��P��.�PRM_�"����HTTP_���H1o (��OcBJ� ��)$���LEyc��d�p � �睱AB_��T@S��S���{�KRLK�HITCOU� À�!퀶������M�SS���v�JQUERY�_FLA!a��B_�WEBSOC�"��HW��a1q�>7�INCPUR�!Ou�ˡ�Č������������IOLN.r 8��R	���$SL2$I�NPUT_PQ$t�ܸP�# ���wSLA�1 sðٿ���s��rNA{IOC�F_AS8Bt$L&��&q�!]�/a�ɳ�@ҳUpHY���lïA�G�UOP5Eu ` X������ā������P������������UQ� M�qqv �l�@;sTAkr��A�TI��.�a�Z0Sն�`PSR�BUZ0ID~0��z���yՏ�!�u�z`w�3��f�G��N��Z0����IRCA��� �x Ĩ��CY�EA{���!���%�R�`�q|�8��DAY_��}�NTVA���i�¦eu��i�SCAepi�CL��������� qy`���ԧb����N_ՀACQ�Ђ�W�rz� O ��������y�G�<]�O! 2y�  ӄ)q{P���P�L�ABzan�Z0t�UN�ISb�PITY0��"ѳ��QIR$6D�|R_URLޏ �$AL10EN��@�� �PH�T�T;_U� �Jt�q} X��t�R��" �0A�D�,J�8FLt@�80�
K�3
�UJR.	5~ ���F|@1w��FgwD��$J�72�O!�$J8B�	7�@\��7s�� 8�	�APHI�@Q��Df@J�7J8�
L_K�E��  �K���LM��  �<��XRK����WATCH_VA�!�pp��FIELDb��y�P&��� �0bpaVyp�ֆCT��E��B`�LG��߁� !��LG_SIZ���@�3@X�O��FD�I� �,Q��]P��� �J&3@J&O�J&�J&�]PJ&�q�E`1_CAM^c�!{@�*h1F���'�$��(�#r��&3@�&O��&��'I�(�(,P�&]P��&�RSI�`  �(/@LN��B�����@{A�g1���K�u1��L~3t2DAU�5EAS�������2�0GH��lQ[�B�OOܑ�� Cr�[�IT8��4<`�n�RE(��8SCRX� ڣs�DIm�SG`nG@RGIPR$D/L@�f�քYB��[�S���Z�W7D[��4f�JG=M�GMNCHH�[�FN�FK�G��I�UF�H2p�HFWDv�HHL�ISTP�J�V�H�P�H�0�HRS"3YHJ��Kc�C4tS �f�x�kG�YUJ��D@jG 3yE�{��BG�I�`PO�WZ&ES�"f�DOC���FEXb�TUI�EI/ ��� /!�dDa�CNc�@��p��� 4	��EpANOGfANA[�ā��AIt瑜��DCASZ���c���bO�hEO�gS?��b�hS�hNHIGN�����A��(��dDE��pTLAL�q��|A��*Є���T�"$���}�h�Ԫ�SA�������ʰ��Z�� �P1
�u2�u3�q���R�`�*І ���V��c ��5�z�x�6��P�6��.�ST��R�0Y���`Q� �$E_�C_�� I�n���8��T)ч Lo��π瀖�x������_�E�NS�_��tD_ �L���X���@���MCh2� =���CLDP��TRQLI��D�2�FLGZ�2�3�f�b��Duf�`�LDf�P�f�ORGjQy�~�(RESERV���Ŕ��Ŕ� #�3�� � 	O�jUA�Ff�SVX0D�R	����'�RCLMC�5�şןG���'�pM�ՠJ�/�3$DEBUGMAS�ÐS�D�"��T�`p�E�� TZ�
�MFR�Q��� � ~�HRS_RU���ځ�A)��UFR3EQ� J�$``�OVERh����v�|P�AEFI���%������ӡ�� \ ��$U���?����P)S�p7 	�C�06��BҒ�G�U�Н�?�( 	"MISC�i� dq1�RQ�5		TBB@�� 1��aa�AX9�!|	�"�EXCES��c۳M��.����9���ܲSC� O� H���_G�@��,��� �2��K��a�|��B@��B_��FLIC��B@QoUIRExSMO��yO��d��ML܀M��� 
��19����5�`pMND�1e�/�o2f2�x��D�#�4INAUT(A�4RSM� ��p�NZ�b!�S^�`0e�PwSTL.� 4��7LOC�RI1P�;EX��ANG�b��n��ODAե��1p�x MF�% 7�+�ۂ|@�e�c0��gSUPᅠqFX/ �IGG�1 � ���ۃb!Cۃ�Vۄ ��V�P���R���R���`���SD�w��TIjȯ��b!M ��� Mt-�MD*��)8��`C�L�@�H�C�GDIA�D�2 W]APC��q��C�D�3)3�qOh�/� a�CU�V����"��OPA_��.� �`t �7㉠f��
 B��P��>P���P���KE�RR�#-$B8�����ND2N�N�D2_TX�XT�RA�cp`��9�L�O�0/�_��	�i2����k��RR2൜� �-��1A$� d�$CALI��c%Gt�a�2�pRIN�!��<$R� SW0�S� `�ABC>�D�_JV ��� 7�_Ju3K
E1SP�$��� PEl3k����� �J`��撚�OiqIM`�ŲCSKPS��� �c�	J�1ŲQ�%�%'�_AZ#��=!�ELNq�N�OCMaP�Ʊ��z0RT���h#�1����1ћ�(o`�*Z�$SM�GMP�n�JG�S�CLB���SPH_@�`Ű+0�#\ � � ORTER��`R� _�`�*�AP@�G�Ų4DIS!�"2[3U�DF�p<1�LWB8VELD�IqN�Z`e0_BL�`��m4���J]4r7�7��4�pIN� �������5QB��
�1��_̰ ��5�2#5l���4z�936ٰDH�B�r ����p$V0� ���#oa$� �l���$\���ൡH �$B�ELN ��!_ACCEs1 �H`��@OIRC_06����NT��/�$PSB�7�L�p��DL� �0�G3�`�F;�I�GD�C�G3�B��E�_�q�PB-P3Q����A_M�G��DDPQ2��FW����ClU�C�BaX�DE�[PPABN6�GRO� EECR�q �_D�!�q�����A�p?$USE_� �c]P�CTR�dY�P�b@"� ��YN߰A a`f�Z�aM����ĵbJPO_0�AGdINC���RpT�ig�.�ENC0L񦲰�A�B��@IN7�I0�B�e��$NT]3�5NT23_@2���cCLOQ0���`-�IP� ���fF0����� ���e��C�0�fMOSI�UQ����3Q�ŲPERCH  s+�2 ]w�hs��rn���@c'["e
P2P�A�B�uL�T�����e��8z�vvTRK�%ʁAY��s��,��r;��0��n&��wbȠMOM��»������S��G��C�R� DU��(RS_BCKLSH_C�r����<v ,�"c��݃�b�1a%CLALM�d��m�@�CHK��NGLRTY��5�d�����_Z�1t_U	M��l�C��^Q�!��n��LMTh_L��V#��j�E��Ð�� ���E���H}���r�&�xPCnq�xH���TUl�CMCv^PbWCN_�Nuc��SFtA�yVb�g��!8��r��<�CATs�SHZ��bT�f]�����f��A�	� QPP�As�gb_Pr�V�_ �� 3�Qp�C�U�F��JG>�X�I�K0OG|V�2TORQU�P �/sL��P��Gr1�P��_W��,��!QAٴPBCصHCصI�I�IHCF$�˱�-��ZPVC�@0����N��1T�RPh�$!Z�JRaKT̙ƴ�DB� �M���M��_DLBA�rGRVߴ��BC��HC��H_����@��COS�p �LN��6�W�=�B@8ٵ @8�
�t�b�(���Z1�Gv��MY?Ѳ��=|'���THET0uNK23HC��<C@�[CB�CB<CC� AS�'�
�5�BC5���SBBCS��GT	S��QCo/��'�x�'��q�$DUC�@�w���t5��5Q�qY_��NE��AAKS�z)!8 @��A����'����LPH����e��SW�o�b� o�q���֙�����EV@�V5�2@X�Vg�UVt�V��V��V��V��V��H@�Y�_PW�ܡvt�H��H��UH��H��H��O1��O@�O�	V�Og�O�t�O��O��O��O
��O��F��"�~b���3�SPBALA�NCE_�ѮLE6j�H_��SP�1S���b��q�PFUL�C�"�"q��:1=�|!UTO_>�F��T1T2B)�B2N %��B�`b$�!f� ��(�B}C��T�pO50�A>ɰINSEG�B q�REV�& p�aDI�F��91��'321�	�OB�!	��Ó��2���`0���LCHgWAR�R7BAB%�~��$MECH+���9a?1T�AX9�P��X6�#B7 � 
pY2��{A�eROBQp�CR�r�5M� ��CyA_A�T �� x $WEgIGH6`�$1�d�3X�I6a�`IF�QNjPLAG'b�S'bܲ 'bBILEOD�o�#p�2ST�@�2P�!	��0`@Ơ�1�0���0
�`yB(aA� � 2�.t�6DEB�U�3L�@<B��M'MY9�E� N��D��$D�Axq$��@S���  ��DO_�@A�1� <�0VFL U�(a�IB&B@N�c�H_p�(`�CBO� �/� %��T�`�a⊑T�!~D�@TICYK�30T1�@%NS���WPNQp1 �CQpR�Ԁ(a!2iU!2uU�@P�ROMP6cE� $IR��&aL�8�R�p�RMAI��aa48b�U_@�S� tB�:`R��COD[CsFU.`�6ID_pp�e� �R�G_SU;FF
� Ca�QdRDOlW� mU @lVGRC!2Id�S Ud!2`e!2le��Id�D�e@��0H� _FIvZA9�cORD&A3 �0�B36��b|&a�@$ZDTe� 	
CA�E�4{ *�!L_NAQ�WPriUDEF_I )xr�V5tuU-BhV7D`hVasuUou�VIS��@���A��hT�suS3tD���D4l���7BD5 (���t[CD��O��BLOCKE�Cci_`{_�W�qIbC`UMHe rIdasIdouId�rUb K�TeDsUdtUb5F�� �q`c,0B�`er`eas `c���EhPP� �t,P�q��@W*�)� �	 �TE���D� ALOOMB_C�^�0�2wVIS!�ITY�2�AS�O'CA_FR1I2#��� SI�q��B�RTP��_P��3tC
�2W��W��������9_��jaEAS�3jb@d������p�R��4���5��6�3ORMU�LA_I��G�	w� h �N7��ECOEFF_O ;Q� ��;Qr�G��3S�0�BCA �O�C�CAGR�� � �� $ �u"�BX+PTM�� �AR(�,%��CER� T	�tn�`�  +"LLkd:�pS�_SV�tw�$L��`���v��`�� ��SETU�sMEA�P(`F��0�CA�b�0� � ���0 �@o��Q2��q�rWP�q�	�tբܑubÕQ��p�q�p+���� ��PREC�a� ? �MSK_���� P�11_USER^!�"}�0��}�^!VEL"�}�0ȥ�!1I�`J �M�TQCFGs�� � YP� OG2NGORE�0P���0~��� 4 ݳ8B7�2H1XYZ�cJ!�o yC�1��_ERR��1� �I�Q�P�ۣ@�aAi����@B�UFINDX� �;�MOR� H�0CU@�QH1����Q�a���"�a�${0��~q����;���G� � $SIj����P��!��VO����0O�BJE���ADJ1U�B�� �AY�p5��D.�OU�`Վ�\'a�b=��T� p]��\��BDIRa��i�� ��"�0DYNH쒣2��T6 �R���,P&@��OPWO}R�� �,�@�SYSBU �SCOP��cҎ���U��b� P ����PA�����C2�OP^`U��!��!XB�AI�IMAGS��0U�7B3IM��o�IN��@�~n�RGOVRD��	��K�PM�m�0� P߀�s��H2L�B=�|� �PMC_E�`cъANM��A�B11�B�@��SL�t��� ��0OVSL:�&S�DEX�q}p"/2G2� ��_��G �`��G�`Qfa�B�C�0p�%�c��/_ZER�����s�� @вb5O&`RI��s0
��P��	��qPL�Ĵ�  $FRE�E��E�������!�Ls����T<D0;@ATUS㰤AGC_T��r�UB� _H��s�A4�`t��� D�AI�2RL���a2S�an S���X�EY������ �0XUP��p�qCPX�PF�D3��^� �PG�Ÿ��$SUBGb5���G�JMPWAIqT�V_%LOW�8BQ��@CVF�QZP�G2b!Rz���U3CC� R��MR�'IGN�R_PL�DBTeB;@P�qH1BW�Pd�$��UP�%IG0�z�PIG3TNLN�&"2R�����N�P)�PEED�8HA�DOW;@�����E�7S4F1!4pSPD.s�� L�0AV�5ps0�3UN�0"+02!R��LY�`� �Q���P��v1��G�$��M�P�@L\+�NPA�T�2�xD��PIP%w0�>��ARSIZ�T���c|q�Om`�h�A�TT���"\�B$�M�EM�B�A>C�3UX���e�PL`�ļ� $���SWIT�CHZ"�AW��ASr�B�BLLBv1��� $BArZ�D�s�BAM� h���I��@J50�����B6�F�A_KN�OW�3R��U!�A�D�H۠~0D��5YPAYLOA鱱�SS�_s�\W��\WZYSL�A�mpLCL_�� !���R�A����T���VF�YC�K��Z貓T��I�XR�M��W_ҬTB���JL)a_J�Q����AND^�9�8d�R�Q����PL�@AL_ ��@~0���A��k�C"�DXSE!��sJ3M`af� T���PDCK��r�C}OŰ_ALPHqc��cBE��W�qo�l ��Т�!�� � ��40R_D_1YZ2�TDŰAR�4x!uxEv0s��TIA4_yu5_y6"�MOM��@ks�sxs�s�s��Bv �ADks�vxs�v�sPUB��R�t�uxs�u��r�Fp��� L$PI�1s��^WP.��xY.�I:�IH�IV�<p}Q7��!�� !��b�ӆ��73HIG�C73w%p4І p4w%� z�І�߈�!x!w%SAMP����B�ЇC�w%�@>c 5�q���7 �Ҁ�  ��p0"p��0p�������hp���	���IN ќ�&�ؘ��ϔw"ښ����:�GAMM�ƕS[%�$GE�T��o��D�d��
�ϡIB��2I0�$HI�_��sЩү��E�м�A��٠ʦLW�����٩�ʦ�b贆0caC�%CHKh��� 	��nI_%� ����\bxΑ�����s����v���c ��$�h 1���I>� RCH_D��'� �$)�LE��������hذ�0MSW�FL�$M�`SCRF
(75_����3�� dƧ���kp��x�p0�����SVv1�P���v�Kǿ�	���S_�SA�A�����NO�`C���d���� d_v_\�J�:ۂ�+R��w�0sD<�4���40�� zʴ�ʈ��چ�1��� �ՕәS�Ak0L���� � ��YL,�a������-��� -���b��9�az�HK����W�{����py�Ȳ�M� ��P��`a�$ 7��"r�M���� � �$���$W���ANG]�Q���d���d@���d��d� נNPP���C��ϐX�0O�c�ΑZq��� �� -�<�OM��"���1�C�U�g�bpCON���0}C�a_�B� |�a�����y7xs7 �s��dzdO~z�A��� J���Ǡ �PP A�PMO�N_QUG� �{ 8�0QCOU��nǀQTH� HO&�n� HYSD@ES�BF� UE� ��@O5$�  �@P�৥���RUNZY�0 O��� � POP+�%����2ROGRA(��x@:�2�Ov+�IT�xINFO��� �A_��8�ȫ�OI�� =(ʰSLEQ�����b�S_ED�d � � ���r�KԙQI#��EȠNU�'(AUT��%COPY�Q��8,����M��NB F+U�PRkUT� I"NF2U�B$G0�$Xa�PRGADJ!�fBX_��2$�0(�&~��&W�(P�(���&73� �NH`_C�YC���RGN�SD���LG�Ob��`NYQ_FREQ�rW����^1RD)L�P:BV0�!�s���CRE���c��IFH�jNAK��%�4_G�STA�TU å�MAI�LI�S&@V��ǀL�AST�1�a04EL�EM:1� �EaN�AB�0EASI &A��v�n�?�B���GF�����I���U2`���� �|BAB�C	PRS�LV	A�Fa��I���qU����JP�'c�FRMS_TRvCΑ��Ci�����A�D E���& 	SB 2�  �V��9V(b8WR���RNTdW&�
�DO`�P�W}�
�22PR �z;0��GRID}��BARS��TY�'C��O�p!� _�4!� �R�T�Oo�74� � |� PORXc�.	bSRV�0)(d fDI��T!pAaTd���^g��^g4\i[�^g6J\i7\i8@aFj��:1�$VALAU�C��9D��F65�� !"E��lb�S�1��_@AN����b�1R c17ATO�TALH��qCsPW�K3I�QYtREGENWzlr�X�H@c5v� TR�C�WqC_S���wlp\CV�!p���u���1GRE�3��P�6B+.  sV_�H�PDA���p�S�_Y�i�o6SV�A�R��2� �"IG_SE�3�p b�5�_/�tC_�V$C�MP���DE�M���Ie�Z��^��zF�HANC�O� p&Q$E�2���INT?`iq��yF%�MASK=�.�@OVR�P� �P ��1Α�W!��T� 4� �_XF�{�V��PSLGV�:1� @K��p5a���Ap�JpSh��4��U0>�!����TEa��`G���`�U�Jd�<��3IL_M~4���p� TQ� �����@-�\�V4�CB�Ph{�4AL�Mc�V1b��V1p�2�2p�3*�3p�4�4p�����p:����p��j�|�IN�VIB��<�)�T��0�2,�28�3,�38�4,�48� hR�ґ��� �T �$MC_F�  ����L����ׅ7pMb8�I׃���S ( ���n�KEEP__HNADD��!�$�@��C��0��Q��?��O��| ��p�p�܇�REM'�IqbL�c�h�U��4e�HPWD w �SBM�~�PCOLLAB���p��5q�2�IT�50`�w"NO��FC�AL��� ,��FL�A$SSYN���M� Cq���XpUP_DLYz!�DELA?дJq�2Y� AD����QQSKIP��� �`-O;�NT�]�i�P_-V�� ^U�*����q���q�� u`�ڂ`�ڏ`�ڜ`��Щ`�ڶ`��9�!�J�2R0� �L�EX�@TX3N�7AN� ��N�}� RDC���� ���Rz�T#OR� ���R�1��x���;TRGEA�r8h@��RFLG�^��5�ER���SPC��1UM_N��2/TH2N�Q�A�� 1� ��A��Q62 � D�Kш��@2_PC�3]�S���1_0L10_C}2��2���7 �� $b�  ���	ViR����0�� �\Ub����m8rj��C1��*=��ID� Gy�XUVL1a�1n��� ;10c�_DS�����<��P�11!� �l�����#C��ATE��$�Q���f���;T�3�HO�ME�� f2n�t������3n��'9K,0f4n�n������ f5n���/!/3/E/
�6n�h/z/�/�/(�/�/�7n��/�/@	??-???c�f8n��b?t?�?�?�?�? �fS���!�  �Ag�p��;�zc�Ed� TC�tD:vtCIOꑔIIt@f�O��_OP�E�C4rlC��POWE�� ^@�l�q�`5�5s ����B$DSB��GNA��3s:�C��b0��S232zE� ����5���ICE;US=sSPE(��a�PARIT �2qO�PB���bFLOWFO�TR9@?rt�UX��CUuP���aUXT���a�ERFAC�ZTT�U.p �2PCHa� t�఩�_`Py���$L ��pOM8���A��8�𥀯�UPDư��f�qPTU@��EX��8#hc�EFA8�����BSP�P�a��|�`�7$USA�X��9��EX�PI��$(`�pY�eR_$�q�`mQ�fWR�OI�D���f��FFRI�END��L�$U�FRAMc�pTO;OLvMYH��r�LENGTH_V�TE�dI�;s��$Z pJxUFIN�V_^ ��_ARGuI%���ITI��bBwX�Sw�vG2�gG1�aꀎc�r�w�_r�O_XP��L�+q4���N�Sc��Cp�Pr�q��G���Rǁ󐒧�XQ؂��h�U���U�������PUd�X nm`E_MG`CT�c�H��h���U�dScG��W�`ć��لD]и@KȅJӂй�������$-� 2!���an �i1�h�`U2�k2=�3�k3�j -����iK���F�`l�P�`x�|�NtV�uV�ТPqC,��r�P��� �V������R��pr�.���E9�<�Os�)E$A��T�P!Rh�U�k�ǓS��P����Sb;Q� ! �ႃ"��K��"����S`�p�p��
 ��$$C��S�������9�9� }ؠVERSI�`����i���I#PP��AA�VM_�a2 �� 0  �5�V�b��S��� ��	 ������9� �����ζ����ϧ��0R�d�l�0�BS^ r�1�� <@ϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� ����������'�9� K�]�o����������� ������#5GY�k}����|�C]C`XLM�@�����  d�IaN����qEX?��2_`=� �9��0�IOCipq ��PZXQ��{�IO'PV 1]=�P $-��ұ0�!̺ �?���  ��//%/7/I/[/ m//�/�/�/�/�/�/ �/?!?3?E?W?i?{? �?�?�?�?�?�?�?O O/OAOSOeOwO�O�O �O�O�O�O�O__+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9oKo ]ooo�o�o�o�o�o�o �o�o#5GYk }������� ��1�C�U�g�y��� ������ӏ���	�� -�?�Q�c�u������� ��ϟ����)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{���ϟϱ���� LAR�MRECOV �I��LMD/G �����_IF  ���p߂ߔߦߴ��^���������, 
 �G���� m�����$_��� ����� �2�D�V�h���NGTOL  �I 	 A �  ����� PPI�NFO %�� $������  1�I
�8r \������� &W�p�Rdv �������/�/*/x�PPLIC�ATION ?�����LR Han�dlingToo�l y" 
V9.10P/25���5'
88340�z#�*F0�!�/13�1y#�,�/�"7D�F1� 5,y#Non}e5+FRA5/� 6�-B&_A�CTIVE��  �[#��  X3UT/OMODb0)���U5CHGAPON�L�? �3OUP�LED 1M��� �0�?�?�?O;CUREQ 1	M�W  TILL�	XOiE_ ~D�;B�m%MD�H6E�2cJHTOTHKYwO��D\COUO_�O7O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_oo#o 5oGoYoko}o�o�o�o �o�o�o1C Ugy����� ��	��-�?�Q�c� u�����󏽏Ϗ��� ��)�;�M�_�q��� ���˟ݟ���� %�7�I�[�m����� ��ǯٯ�����!�3� E�W�i�{���翱�ÿ տ�����/�A�S� e�wω��ϭϿ����� ����+�=�O�a�s� ���ߩ߻����������'�9�K�CETO��d?X2DO_C�LEAN�?V4��N�M  �� �O*�<�N�`�r�ND?SPDRYR��U5HI�0�@����� &8J\n�p���R8MAXI  ��|�~A�7�X���!��2�!X2PLUGGp�0���3t5PRC��B�����.�O3����SEGF�0Kz�������//&/^�LAP����Cz/�/�/�/ �/�/�/�/
??.?@?|R?�3TOTAL�|�3USENU���; ��?~B@R�GDISPMMCʚ�AC��@@$���4O�����3�_STRING �1
�;
��M�0ST:
)A_�ITEM13F  nT=OOaOsO�O�O�O �O�O�O�O__'_9_�K_]_o_�_�_�_�I/O SIGN�AL-ETry�out Mode�4EInp�PSimulated8A�Out�\O�VERR�� = �1007BIn �cycl�U8AP�rog Abor�c8A�TStat�us6C	Hear�tbeat2GM?H Faulug~cAler�i�_�o�o �o�o�o $6H ��/K��AOK �������� )�;�M�_�q�������p��ˏݏ_WOR� /K���=�O�a�s� ��������͟ߟ�� �'�9�K�]�o�����PO-Kia��-��� ܯ� ��$�6�H�Z� l�~�������ƿؿ����� �2ϴ�DEV ��]�ЯJτϖϨϺ� ��������&�8�J� \�n߀ߒߤ߶�����PALTu}�-� ��)�;�M�_�q��� �����������%��7�I�[�m���GRI � /K���������� '9K]o� ����������0Ru}I��#q �������/ /%/7/I/[/m//�/x�/�/7PREG� � a�/?'?9?K?]? o?�?�?�?�?�?�?�?��?O#O5OGOYO�]��$ARG_�D �?	����A��  w	$�V	[�H�]�G��W�I�@SB�N_CONFIG(�P�K�Q�RQ�A�CII_SAVE�  �TQS�@T�CELLSETU�P �J%  ?OME_IO�]�\%MOV_HVPi_o_REPL�_�JUTOBACKAQ��IQFRwA:\�+ �_,�&P'`T`�'h�� k
P �18/02/�09 11:06:04�&�H�-{o0�o�o�o�\���o@%7I[�&��o ������n� �+�=�O�a�s���� ����͏ߏ�|��'��9�K�]�o���X� � �Q_�S_\AT�BCKCTL.TM����ҟ�����[INI�AeV�S?MESSAG!P/��Q�@SQD�ODE�_D[P$VUb�Ox_�q��SPAUS͠� !��K ,,		��@�Eѯߧ ů������Y�C� }�g�y�����׿��ӿ��������TSK�  ��o��PUgPDTh�-�d~��~�XWZD_ENqB-��J��STA,���A~ŎAXIS�@U�NT 2�EQ�P� 	D�
V����5�� �$z�9� ֘Y�*��  "�ASXjE�!*�=��O�����@�~� ��$ ~�9Bv 2�r,�RU�%2h6߸�߉F��METK2�4�-S P��B��>B���C
�AH>l�ZB��M�B�K��@�@4?6��?��]>]0�?Lc@@�����SCRDCFG �1�E�Q 	�)UR�߆��� ������o�*Q%Ys� 0�B�T�f�x������ �������,�����G�QGR��r����k��NA�P�K	��Th_ED+�1�V�� 
 �%{-��EDT-Y��Z�M�
TzP-(�S��*�B�otV���  ��u2 ~�[\���'�/ Yk/�w3J/� �/��s/�/%/7/�/[/w4?�/c?�/��??�?�/?�?'?w5 �?R?/Ov?�OvO�?�?eO�?w6�OO�O BO��OB_�O�O1_�Ow7z_�O�__��_@oU_g_�_�_w8Fo��o��oo�o!o3o�oWow9�o_�o��;��o�o�#wCR}�_*�<� �]�p���_��k ~� NO_DELw��GE_UNUS�Eu�IGALL�OW 1�	 �  (*SY�STEM+�	$SERV_GR���*���REG3�$8U�Q�*�NUMX�}��k�PMUրQ��LAY��Q�?PMPAL,����CYC10��ʞx�����ULSU��0l�̒��5�L�?��BOXORI\�C�UR_,�k�PM�CNV��,�1�0����T4DLI���%�G�	*PRO�GRA2�PG�_MI�����AL(¥����B�*��$FLUI_R�ESUЗX�b�����������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ����������H�k LA�L_OUT ��T�WD_AB�ORѐ��jO�IT�R_RTN  �st��O�NONS�TO� z� b�CE_RIA_I���z������F?CFG �
���s}��_PA9�G�P 1�����Q>�P�b�!�C��p����z�C�Ce ��(����C8��e@��H�� CX��U`��h��p��x}�U������������	su?����HE��ONFI���Y�3G_Pr�1�� ��ă�} �������3�KPAUSI�1`�� ���C` 1oU���� ���/5//Y/k/�Q/�/Mo�NFOw 1`�� � 	-��/�p�� ��Bv�ſ��X��n²�C~�������	���	�(>B��hC3���9!C2���1��@�D�"(>�N���a�3�]���2����O�����sw�COLLEWCT_���&A���~7EN z���2nW1NDE�3�7�eヂ1234?567890�7~r`D����?�6ss
 ���q)9O^OD�8OJO �OE�|O�O�O�O�O�O /_�O__w_B_T_f_ �_�_�_�_o�_�_�_ Ooo,o>o�oboto�o��o�o�6B�2�;� �=�2IO  �9�1yxy�as�l�/wTR�2!}��� Jy
�o�~> �">}�z���9_MO5Rr#
� �'	X� �!X�p�^����������1� �q$?�,C?$,,��UpK�Tq�Jr��P[2&�?"� +�a�s�����
R���t7���u�y���5����s ���9P�DB/�(7��dc?pmidbg�]�Lv o�:��nD�pI�|��m�  ��n1G�毱��ï��l.�����mg�x�C�Ůfg����-ſ>�`ud1:����z'�DEF '�y(Is)��c�b?uf.txt�g�\�%�_MC8�)7�"!sd�ō�7�*���������|�Cz  B�3A� D��C����C-y�CZ��Џ����-E�d�1E���E�9KD���E�;�#��-G����G�?kGW6��F�NGWeG��|ɰ�Vq���,|��t7ARUpH b�H �H ɐ�t
��� ќ@� Da  D� � E	� D�@� ���-F| F�p F"� G�=�fF��G�'i;�>�G�g� GK  H��<=H�&H�yMc��  >�33  `C/b��n)���5YT�䨂��A�|�=L��<#� �Vq�����ξ��RSMOFS�T %8ʝ/�&P�_T1��DE -3����q��Tq�;������?����<�;��EKST2�+8�PR�2�.a?����C4���|��Up��������mC��B���C�����H�Up:d�� ���T_2�PRO'G ���%x�V�$INUSER � �5($KEY�_TBL  ��"�	
��� !"#$%&'�()*+,-./��7:;<=>?@�ABC2�GHIJ�KLMNOPQR�STUVWXYZ�[\]^_`ab�cdefghij�klmnopqr�stuvwxyz�{|}~����������������������������������������������������������������������������0��͓���������������������������������耇���������������������9�q* LCKt��<&t STAT����_AUTO_DOr�6���IND�4��}1R���T27/�STO@/� �TRL, LETE��7~*_SCRE�EN ?��kcsc�2Uo MMENU 1/.� <ED?[ �/?J?ճ'?M?�?]? o?�?�?�?�?�?�?O :OO#OpOGOYO�O}O �O�O�O�O�O$_�O_ Z_1_C_i_�_y_�_�_ �_�_o�_�_oVo-o ?o�ocouo�o�o�o�o 
�o�o@)vM _������� *���9�r�I�[��� ���ޏ��Ǐ�&��� �\�3�E���i�{����ڟ��ß�Ϲ�#_M�ANUALs/�!DwBCO RIG�'|�/�_ERRL2 0��a�N������ǯ P�NUMLQI;�Z!v�d��
P��PXWORK 11����'�9�K�]�|o��DBTB_�!G 2��ç�����DB_AWA�YX�a�GCP r��=E�ö_AL;��òT�Yr �%��I��_r� 13#� , 
�T��B�ϖ��_M I��Ѽ@|����ONTIM�'��������
��$�MOTNEN���z$�RECOR�D 19�� �<�ψ�G�O�O�=� ��Ҳ{ߍߟ߱�Hع� ��O��s�(�:�L��� �߂��ߦ��������  ���$���H���l�~� �������5���Y�  2D��h����� ����U
y �Rdv��� �?�//*/�N/ 9/G/�/��/�/�/;/ �/�/q/&?�/J?\?n?�?}?�??�?7?����OO�?9O$O�? oO�?�O�O�O&O�O�O \O_�O5_G_Y_�OZ�òTOLEREN�CдB��ްL���P�CSS_CNSTCY 2:�%���i_���_�_ �_oo'o9oKoaooo �o�o�o�o�o�o�o�o�#�TDEVIC�E 2;�[  ��vu���������*��ϭSHN?DGD <�[��Cz|{�TLS 2=]}<�����Џ�����>��RPARAM >0� |���}�SLAVE �?]�I�_CFG� @J�*�d�MC:\�PL%0?4d.CSV)�頱cџ�RA ��C	H�o�o�*��F��w�76��1s�a��1�JP��3|����r�_CRC_?OUT A]}��~.�_NOCOD~��B0���SGN �C&��&j���21-APR�-21 01:2�4�*�09-�FEB-18 1�1:06��v LIX�v�r�*��s�Iu5�M���Þ���������VERSI�ON -�V4.2.10���EFLOGIC {1D�[ 	�8�+�ɘ�!��PR?OG_ENB�e��A�ULS�� d���_ACCLIM^��������WRSTJNT���*��MOJ������INIT EؼZ&�*� ��OP�Ty� ?	����
� 	R575�*�+�740�61�7R1�5�[�1U�21���8���TO  �݉����V��DKEX��d��Hp��?PATH ۦ�A\��9�K�[H�CP_CLNTI�D ?Ѷ�� ��? ��RIAG_GRP 2J��� Q 	� @K�@�G�?���?l?��>���� ���Q ����ᴝP)�>�?�b�?PT��i�^?�Vm?�Sݘ��f4�03 6789012345{������� ��s��@�nȴ@i�#@�d�/@_�w@�Z~�@U/@�O�@I��@�D(����@�b��p����PA�PY�P�B4��jp���ط�
��1��-�@)hs@$���@ bN@��@�����@�D@+ ����������	 ���R��@N@�I�@D�@�>�y@9��@�4� .v�@(��@"�\Pbt���L�@G�l�@BJ@<�z�@6��0�`�@*� $N�@��� |$=q@����F@|�@�33@�R@�-?���?��`?�+h�z����Y"J��-@&�@�N���!?�??� ��/ /*/</�-�/?�/ &?8?�/?Z?�?^?�? �?@?R?�?�?O�?4O FO�?VO����9��Q�i @��V�AY�����?�z��A��5AF�A4���@��L4Ry��A��@�p� R�Q�R-PP���@�� ��Ah��=�H�9=Ƨ�=ߺ^5=�>P���>���=��,d_�,P� ����C��<(�U�\� 4����_�-���A@��?��pO �_xM�_o0o�ȡT<o fo ovo�o~o�o�o|I�>��y�b�R�=���=��z�q���G�G��� � ��!�!�NUt�@�T��V��u�B�� B��B��B%������~'���up���q�q6|�\�&����g���)PB3pBj�B A�@�"����m���<�� � ��e<�)_N�3���?���6_�67<U�6[�����C	���	(@B���]�l���r�ݏȏD��x�"������C3��9 O��C2��@Cҿ ��q�쏕�������ݟ�ȟN�PB>�)�'<�ٗ����?�ܿ�*xM��=���CT_CON?FIG K�m��eg7Ų�STBF_TTS�ǁ
YɈ�Ȱ���������MAU��N���M_SW_CF\�L���  ���OCVI�EW��M������A�S�e�w����� ��/�Ŀֿ����� ��B�T�f�xϊϜ�+� ����������,߻� P�b�t߆ߘߪ�9��� ������(��L�^� p�����G�����  ��$�6���Z�l�~��������D�RC�N(E��!P�����!�E4iX���SB�L_FAULT �O����GPM�SK���P�TDI�AG P`��q�o��o�UD�1: 6789012345t�n���P*�Sew� ������// +/=/O/a/s/2����R
B�/�TRECP�
?) �+A>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^O�/�/�/�O��UMP_OPTIcON����ATR�t���	�EPME����OY_TEMP  È�3B��5P��TUNI�͠��5QܦYN_B�RK Q��EDITOR�A�A_��R_� ENT 1�R��  ,&�PROG ANIE2 M�Q�_�D��PICK�_o &DROP�_�3o`
ZEROW�#o`o&}�os��to�o�o�o�o�o �o/SeL�p ������� � =�$�a�H�p���~������ߏ�؏����PMGDI_STAHU�$�5Q}UNC;�1S� �dO��v��N
�Nd�Oݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W��En��������� ʑ��ؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@ߺ� g�q߃ߕߧ������� ����%�7�I�[�m� ������������ �!�3�E�_�i�{��� ������������ /ASew��� ����+= W�Es������ ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?Oak?}? �?E?��?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ G?Y?c_u_�_�_�?�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7Q_[m ��_����� �!�3�E�W�i�{��� ����ÏՏ����� /�IS�e�w������ ��џ�����+�=� O�a�s���������ͯ ߯���'�A�3�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �9�K�U�g�yߋߥ� ����������	��-� ?�Q�c�u����� ����������C�M� _�q����ߧ������� ��%7I[m ������� !;�EWi{�� ������// //A/S/e/w/�/�/�/ �/�/�/�/??3!? O?a?s?��?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O_+?=?G_Y_k_!_ �?�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	#_5_ ?Qcu�_��� �����)�;�M� _�q���������ˏݏ ���-7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����%� /�A�S�e��q����� ��ѿ�����+�=� O�a�sυϗϩϻ��� �������9�K�]� w����ߥ߷������� ���#�5�G�Y�k�}� ������������� '�1�C�U�g��ߋ��� ����������	- ?Qcu���� ���m��);M _y������� �//%/7/I/[/m/ /�/�/�/�/�/�/�/ !?3?E?W?q{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O?�O+_=_ O_i?__�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o __#5G�os_} �������� �1�C�U�g�y����� ����ӏ��o�-� ?�Q�ku��������� ϟ����)�;�M� _�q���������˯ݯ �	��%�7�I�c�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ���������� /�A�[�M�w߉ߛ߭� ����������+�=� O�a�s������� �������'�9�S�e� o��������������� ��#5GYk} �������� 1C]�gy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/I�??)?;?U _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�/�O _!_3_M?W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�O�o+E_ ;as����� ����'�9�K�]��o���������ɏ�o ��$ENETMO�DE 1TFu�  �`��`�e�"��R�ROR_PROG %��%�fe�r��@�TABLE  ��P��ß՟��@�SEV_NUM� �  ��	��@�_AUT�O_ENB  �,��=�_NO� �U��!�� W *�]��]��]�	�]��+\�v������6�FLTR"�4�H�IS��a�/�_A�LM 1V�� e��d]��`+���6�H�Z�l�~�����_\��<�  ��[��"�պ�TCP_V_ER !��!]����$EXTLOGo_REQ֦�-��'�SIZ0�"�ST�KM�K��$�T�OL  �aDz�ޢ�A "�_BWD��������'��ûDI�� WFu��� ��a��ST�EP�������OP�_DOo���FDR_GRP 1X����d 	пm�"�^��n&���c�?��$,�MT� ��$ �����^ӳ����^�B�8 B���!C ��B�"dB\�vB%���� $B`��B���Aб�A�e(A�ŷ ����:�%�^�I��m�����  A,�f�At�>(������`
 M�q�	����ⲉ�������?�*�c���A�@����@�33@%�������@����L�����^�F@ ���E��������L�FZ!D��`�D�� BT���@�����?�  M��6����u��5�Z�f5�ES�����e�����J �9���`�Zy�w�>x�FE�ATURE Y�Fu��&�L�R HandlingTool ���bEngli�sh Dicti�onary�4Dw St� ard���Analog �I/O#,gle� Shift?u�to Softw�are Upda�tedmatic Backup�	��ground �Edit� �Ca�mera:F>C�ommon ca?lib UI���n��Monit�or�tr� Re�liabS�DH�CP��
Data Acquis�~%)iagnos��7?+ocument Viewe"�''ual Che�ck Safet�y��hance�d��
�%s� Fr���xt. DI�O �fiu$�'e�nd� Err L(t"	=�'s9r5� � ���
FCTN /Menu� v##[7�TP InJ0faycq5�GigE�>��5�p Mask� Exc� g�'H�T�0Proxy �Sv�$�6igh-wSpe� Ski���6m � mmuni�c�onsHur�h0J0:/;�2con�nect 2:Hn{cr�0stru$8Ja@e�!� Jt%��KAREL Cmod. L�0ua�8~�CRun-Ti� �Env�HK0el u+�s�S/W�License�#��,0Book(S�ystem)�
M�ACROs,�2/�OffseZUH0� w8/"PMR ��s.M}M@!l�,MechStop�1tQ@Y"Ui2V�Vax� 7�L^odTwitch�_aSh!y.BV�[OptmoLaS�0fi�^aVg0G~Uulti-T�0���	PCM fu�nkG�ia�Ptiz�~h�goV$Regi�Pr@�fri� F��k�f8Num S�el�U�i�  Ad�ju@�n qV1}t�atu�aI�*�R�DM Robot>scove�u�eav`� Freq� AnlyGRe�m�P�!n�u�rS�ervo� �P�S�NPX b�B[SN�0Cli�!�W�Libr(��  ��T:��vo�@th0sGsag~e�� l�5Q&�/I�=��M�ILIB����P OFirmu��Ph3�Acc��TPT9X4/��eln5PǏ����1U��orqu>Timula!�E�u�PPa�A���t!!c&�0ev.���mri� �US?R EVNTğ֐nexcept� ��pn�#ѕ�(@VC"�rBB�XVU 6���G�:�A�S�SC��y�SGE����U�I&Web Pl `vǮ�q0O��0�$�!�?6ZDT AppYlD�
iP0a!��:� Grid�qp�lay=����W�R-�.��h!N��B^P�}200iV4+s�cii�1rLoa9d� �Upl����f@I�Pat�V�y�cS�B�`��� \6R�L��� ۩�5MI 7Dev�@ (�qRx�f�?�gsswo!��_64MB D�RAMM���FRO��Ͼell:�sh��#�c.k �rYp��5�tySs
r7̬r'`.?+�p�!"�=-o� 2�a5p�ort�.�p�r q�-T1 �{]P��ONo m�pc$�v��OL��Sup���Fa�hOPC-UA��l�T �2eϓ�S0�0croa|�s:�����~���uest��uS��e2tex�V��up�1�#��PPx�00�oVirt�!|�sR�stdpnÛ��� SWIMES7T f F0�����������������  MDVpz ������
 I@Rlv�� ����///E/ </N/h/r/�/�/�/�/ �/�/???A?8?J? d?n?�?�?�?�?�?�? O�?O=O4OFO`OjO �O�O�O�O�O�O_�O _9_0_B_\_f_�_�_ �_�_�_�_�_�_o5o ,o>oXobo�o�o�o�o �o�o�o�o1(: T^������ �� �-�$�6�P�Z� ��~�������Ə�� ��)� �2�L�V���z� ����������%� �.�H�R��v����� ��������!��*� D�N�{�r��������� �޿���&�@�J� w�nπϭϤ϶����� ����"�<�F�s�j� |ߩߠ߲�������� ��8�B�o�f�x�� ������������ 4�>�k�b�t������� ������0: g^p����� �	 ,6cZ l������/ �/(/2/_/V/h/�/ �/�/�/�/�/?�/
? $?.?[?R?d?�?�?�? �?�?�?�?�?O O*O WONO`O�O�O�O�O�O �O�O�O__&_S_J_ \_�_�_�_�_�_�_�_ �_�_o"oOoFoXo�o |o�o�o�o�o�o�o�o KBT�x� �������� G�>�P�}�t������� ��������C�:� L�y�p���������� ܟ���?�6�H�u� l�~��������د� ��;�2�D�q�h�z� ������ݿԿ� �
� 7�.�@�m�d�vϣϚ� �����������3�*� <�i�`�rߟߖߨ��� �������/�&�8�e� \�n���������� ����+�"�4�a�X�j� ���������������� '0]Tf�� ������# ,YPb���� ����//(/U/ L/^/�/�/�/�/�/�/ �/�/??$?Q?H?Z? �?~?�?�?�?�?�?�? OO OMODOVO�OzO �O�O�O�O�O�O_
_ _I_@_R__v_�_�_ �_�_�_�_oooEo <oNo{oro�o�o�o�o �o�oA8J wn������ ���=�4�F�s�j��|�����̍  ?H551��⁽2�R782�5�0�J614�AwTUP�545��6�VCAM�C�UIF�28H�N�RE�52;�R6�3�SCH�DO�CV��CSU�8�69�0�EIOuCl�4��R69;��ESET$�:�J7�:�R68�MAS�K�PRXYT�7.�OCO�3$�������37�J6
�5u3��He�LCH��OPLG$�0O�M�HCR �S��MA]Tk�MCS#�0��{55�MDSW�vB�OPB�MPRC�t��s�0�PCMS��5J������s�51�/�51{�0/�PR�S�697�FRD�G�FREQ�MC�N�93�SNByAx�f�SHLB��M
ǀ���2�HT=C#�TMIL􈳖�TPA˖TPTXF<�EL۶����8������J95_�TU�TC�UEV�UE�C�UFRG�VCuC��OǦVIPG�wCSCk�CSGk����I�WEB#�H�TT#�R6v���C�G6�IG�IPGmS\�RCG�DGB��H75/�R7�R�y�R66O�2O�R]6�R55��4��]5��D06�F��CLI3�.�CMS�˖0�#�STY��T�O7�7��t�_�OR�SǦ��M��NO�M˖OL�$���O{PIs�SEND�uL��Sy�ETSs�켐S�CPk�FVR�˖IPNG�Gene�È6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� ��ԟ���
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲����������� 0�B�T�f�x���� ����������,�>� P�b�t����������� ����(:L^�p�����	 � H551���2�
R782��50�	J614��	ATUP54�56�	VCAM��	CUIF28nlNRE�
52[wR63�SCH�	�DOCV�CSU��
8690+E�IOC�4R6=9[ESET<Z�J7ZR68�
M�ASK�	PRXY�|7�
OCOL,3�<X 3�*J6�53�H�,LC�H�*OPLG<0^�*MHCR�*SJ;wMAT�MCS;�0[+55+MDS�W�;�+OP�+MP�R�*��,0PCM{5KX +X0�+[51K51[L0K�PRSK+69�*F{RDkFREQ�
�MCN�
93S�NBA��+SHLEB�JM[��<2�HTC;TMIL���TPA*TPTX\ZEL�JX0�q8
�
J95�wTUT�*UEVK*wUEC�*UFRk�VCC+lOk:VI�PkZCSC�ZCS�G��I�	WEBn;HTT;R6���\CG�kIG�kI�PGS�jRCkZD�G�+H75KR7�:+RYLR66�,2v�*R6�R55k|u4�[5�{D06+�F�|CLI�<JC�MS*�p;STY[kTO�k7���GORSk:x M�L7NOM*OL�;�0��OPI�jSEN�D�
L:kSY�ET�S�j {[CP�F�VR*IPNkZGene��R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&� 8�J�\�n߀ߒߤ߶� ���������"�4�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt�И���� �STD�LANG��	'9 K]o����� ���/#/5/G/Y/ k/}/�/�/�/�/�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	O O-O?OQOcOuO�O�O �O�O�O�O�O__)_�;_M___q_�ZRBT�OPTN�_�_�_|�_�_DPN� oo*o<oNo`oro�o �o�o�o�o�o�o?ted �� >Pbt���� �����(�:�L� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����*�<� N�`�rτϖϨϺ��� ������&�8�J�\� n߀ߒߤ߶������� ���"�4�F�X�j�|� ������������� �0�B�T�f�x����� ����������, >Pbt���� ���(:L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/�/ ? ?2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_ �_�_oo&o8oJo\o no�o�o�o�o�o�o�o �o"4FXj| ��������8�0�B�  �K�i��{�������Í99�ʅ�$FEAT_�ADD ?	��������  	ǈ��,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O��O�O�O�O�O�O�D�EMO Y��   ǈ1]'_ 9_f_]_o_�_�_�_�_ �_�_�_�_,o#o5obo Yoko�o�o�o�o�o�o �o�o(1^Ug �������� $��-�Z�Q�c����� ��Ə��Ϗ�� �� )�V�M�_������� ��˟����%�R� I�[����������ǯ ����!�N�E�W� ��{�������ÿݿ� ���J�A�Sπ�w� �϶ϭϿ������� �F�=�O�|�s߅߲� �߻��������B� 9�K�x�o����� ��������>�5�G� t�k�}����������� ��:1Cpg y����� � 	6-?lcu� ������/2/ )/;/h/_/q/�/�/�/ �/�/�/�/?.?%?7? d?[?m?�?�?�?�?�? �?�?�?*O!O3O`OWO iO�O�O�O�O�O�O�O �O&__/_\_S_e_�_ �_�_�_�_�_�_�_"o o+oXoOoao�o�o�o �o�o�o�o�o' TK]����� �����#�P�G� Y���}���������׏ ����L�C�U��� y�������ܟӟ�� 	��H�?�Q�~�u��� ����دϯ���� D�;�M�z�q������� Կ˿ݿ
���@�7� I�v�m�ϙϣ����� ������<�3�E�r� i�{ߕߟ�������� ���8�/�A�n�e�w� ������������� 4�+�=�j�a�s����� ����������0' 9f]o���� ����,#5b Yk������ ��(//1/^/U/g/ �/�/�/�/�/�/�/�/ $??-?Z?Q?c?}?�? �?�?�?�?�?�? OO )OVOMO_OyO�O�O�O �O�O�O�O__%_R_ I_[_u__�_�_�_�_ �_�_oo!oNoEoWo qo{o�o�o�o�o�o�o JASmw �������� �F�=�O�i�s����� ��֏͏ߏ���B� 9�K�e�o�������ҟ ɟ۟����>�5�G� a�k�������ίůׯ ����:�1�C�]�g� ������ʿ��ӿ ��� 	�6�-�?�Y�cϐχ� ���Ͻ��������2� )�;�U�_ߌ߃ߕ��� ���������.�%�7� Q�[�������� ������*�!�3�M�W� ��{������������� ��&/IS�w �������" +EO|s�� �����//'/ A/K/x/o/�/�/�/�/ �/�/�/??#?=?G? t?k?}?�?�?�?�?�? �?OOO9OCOpOgO yO�O�O�O�O�O�O_ 	__5_?_l_c_u_�_ �_�_�_�_�_ooo 1o;oho_oqo�o�o�o �o�o�o
-7 d[m����� ����)�3�`�W� i�������̏ÏՏ� ���%�/�\�S�e��� ����ȟ��џ����� !�+�X�O�a������� į��ͯ�����'� T�K�]����������� ɿ������#�P�G� Yφ�}Ϗϼϳ�����|���  � +�=�O�a�s߅ߗߩ� ����������'�9� K�]�o������� �������#�5�G�Y� k�}������������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������� ��������'9 K]o����� ���#5GY k}������ �//1/C/U/g/y/ �/�/�/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?OO)O ;OMO_OqO�O�O�O�O��O�O�O_Y  XQ/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoaoso�o �o�o�o�o�o�o '9K]o��� ������#�5� G�Y�k�}�������ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��������ϯ��� �)�;�M�_�q����� ����˿ݿ���%� 7�I�[�m�ϑϣϵ� ���������!�3�E� W�i�{ߍߟ߱����� ������/�A�S�e� w����������� ��+�=�O�a�s��� ������������ '9K]o��� �����#5 GYk}���� ���//1/C/U/ g/y/�/�/�/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?O O)O;OMO_OqO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/ASe w������� ��+�=�O�a�s��� ������͏ߏ��� '�9�K�]�o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O(�O	_QPX3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c� u���������Ͽ�� ��)�;�M�_�qσ� �ϧϹ��������� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ������� '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����������	���$FE�AT_DEMOIoN   ԀK��� �3�INDE�X@�Oш3�IL�ECOMP Z�������N�.�w�SETUPo2 [����?�  N ��t��_AP2BCK �1\��  �)�����%��� ����H����t�� ��'����]����� (���L���p������ 5�����k� ��$�� 1Z��~��C �g��2�V h���?�� u
/�./@/�d/� �/�/)/�/M/�/�/�/ ?�/<?�/I?r??�? %?�?�?[?�??O&O �?JO�?nO�OO�O3O �OWO�O�O�O"_�OF_ X_�O|__�_�_A_�_ e_�_o�_0o�_To�_ ao�oo�o=o�o�oso �o,>�ob�o� �'�K�o��t����P�� 2��*.VR�g��p*j����s�����u�Q�PC��pF'R6:֏���;�ʋT_�_�q� �\����B�,����v*.F�T���q	����x��C�қSTM c��l�w��d����p�iPendant? Panel��қH������该�3�L�ӚGIFV�����l�p)�;�пӚJPGڿ�ϋ�𿭿��T�ˊJS^χ��p�u�2��%
JavaSc�ript��޿CS��ߊ��ϵ� %�Cascadin�g Style ?Sheets7ߩp�
ARGNAME�.DTf��|��\@z�8ߚ��Ի�g���DISP*�ߔߎ����>���0�?���	P�ANEL15��%������ﵯǯu�2 ����������o�z�3;������L�^���z�4��%�������wr�TPEINS�.XML~�:\��PbCusto�m Toolba�r���PASSW�ORDC�~FR�S:\� %�Password ConfigW��4�/�ԝ[U� /qֱ䘯���/�`b_/v���/%J( �/g/y/?'2T/=? H(+?�/�/�?��?�/@U5�?o?�?O'3\? EOH(3O�?O�O���O��?]E�OwO�O_'4 dOM_H(;_�O_�_ �_�OeU�__�_&o� Jo�no���o3o�o Wo�o�o�o"�oFX �o|��A�e ���0��T��M� �����=�ҏ�s�� ��,�>�͏b�񏆟� '���K���o�ٟ��� :�ɟ^�p�����#��� ʯY��}������H� ׯl���e���1�ƿU� ����� ϯ�D�V�� z�	Ϟ�-�?���c��� ����.߽�R���v߈� ߬�;�����q��� *����`��߄��}� ��I���m�����8� ��\�n����!���E� W���{���	F�� j����/�S� ���B��x �+��a�,��$FILE_D�GBCK 1\������� < �)
�SUMMARY.sDG/�]MD::/�z/�Diag� Summary�{/([CONSLO�Gp/S/e!�/�/�!�Console �log�/�\TPA'CCN�/Y?%A?~?��%TP Acc?ountin ?��Y@6:IPKDM�P.ZIP�?�
��?O�%�0Exce�ptionO�*�_\O�bQJO�_�1FR DT F�iles�O�<f MEMCHECKt?��/i/_1Mem�ory Data�_�l�)	FTP�/f_�Oj_W�1mme`TB�D�_�L >I)�ETHERNE�T�_��A�_o�!�Ethernet� 0figura�&O�}QDCSVR�F�_m__�oQ%�]` verif�y all�o�M�.cXeDIFF��ovo�o P%�hdiff�g�A>]`CHG01�o���a5��b- `y2��&�1���gr3������ <�я`�VT�RNDIAG.LAS֏����.�!Q�� Ope>c Lo�g �!nosti�cCW��)V7DEV�DA}O�x����aVisQ�?DeviceX�e�IMG��?����4�z7�ʔImag֟nc�UP{�ESz�~�FRS:\z���O@Update?s List����"�FLEXEV�ENo�%�>��a�� UIF Ev��QU�?�  ,�s�z)
PSRBW�LD.CMj��𦢂���0PS_R?OBOWEL�_�}*�HADOW4���+�D�SSha�dow Chan�g�ODVa��RCMERR<�!�3����S��CFG �ErrorАta�ilk� a�|�B��SGLIB��ЧϹ�N�!Q� S�t?`_�����):�ZDU_��7���nWZDT�adn�z���NOTIbo�߽�R�UNot�ific?b��t��{AGXbGIGE���/�A���]�GigExZ�d��N�A�� -��Q��^������ :�����p���); ��_����$�H �l��7�[ m�� ��V� z/!/�E/�i/� v/�/./�/R/�/�/�/ ?�/A?S?�/w??�? �?<?�?`?�?�?O+O �?OO�?sO�OO�O8O �O�OnO_�O'_9_�O ]_�O�__�_�_F_�_ j_�_o�_5o�_Yoko �_�oo�o�oTo�oxo �oC�og�o� �,�P���� �?�Q��u����(� ��Ϗ^�󏂏�)��� M�܏q������6�˟ ݟl����%���2�[� �������D�ٯh� �����3�¯W�i��� �����@����v�� ��/�A�пe����ϛ� *Ͽ�N����τ�ߨ� =���J�s�ߗ�&߻� ��\��߀��'��K� ��o����4���X� �����#���G�Y��� }������B���f��� ��1��U��b� �>��t	��$FILE_F�RSPRT  ���� ����$MDON�LY 1\8�  
 ��{� �������/ //�S/�w/�//�/ </�/�/r/?�/+?�/ 8?a?�/�??�?�?J? �?n?OO�?9O�?]O oO�?�O"O�OFO�O�O |O_�O5_G_�Ok_�O �_�_0_�_T_�_�_�_�o�_Co�_Poyo"VISBCKV@e*.VD�o�o8`�FR:\�`ION\DATA\�o�Zb8`Visi�on VD file�oo>Pfot ^o�'��]�� �(��L��p��� ��5�ʏ܏�� ���$� ��5�Z��~������ C�؟g�������2��� V�h�#������?��� �u�
���.�@�ϯd��󯈿�)���LU�I_CONFIG7 ]8�aɻ� $ ��[{ 8 �2�D�V�h�zψ��|x���������� ��
ܠ�-�?�Q�c�u� ߆߽߫������ߊ� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi ����� �~/ASe ������h� //+/=/O/�s/�/ �/�/�/�/d/�/?? '?9?K?�/o?�?�?�? �?�?`?�?�?O#O5O GO�?kO}O�O�O�O�O \O�O�O__1_C_�O g_y_�_�_�_�_X_�_ �_	oo-o�_>ocouo �o�o�oBo�o�o�o )�oM_q�� �>�����%� �I�[�m������:� Ǐُ����!���E� W�i�{�����6�ß՟ �������A�S�e� w��� �����ѯ��� ���+�=�O�a�s��� �����Ϳ߿�Ϛ� '�9�K�]�oρ�ϥ� ���������ϖ�#�5� G�Y�k�}�ߡ߳��� �����ߎ��1�C�U�(g�y�	���x�����$FLUI_D�ATA ^���������RESULT� 2_���� ��T�/wi�zard/gui�ded/step�s/Expert ��"�4�F�X�j�|��������������C�ontinue �with G��ance��1CU gy������� ��-����0 ������6$���ps�o �������� /#/5/���\/n/�/ �/�/�/�/�/�/�/?�"?4?F>$(:Jrip�X�?�? �?�?OO*O<ONO`O rO�OC/�O�O�O�O�O __&_8_J_\_n_�_@�_Q?c?�_�?EJ��TimeUS/DST�_"o4oFoXo jo|o�o�o�o�o�o��?Enabl
 .@Rdv��P������ `�_��_�_f24o r���������̏ޏ�� ��&��o�o\�n��� ������ȟڟ���� "�4����)�;�M�zon
`7�ʯܯ�  ��$�6�H�Z�l�~����EST Ea��rn Stand������ӿ���	� �-�?�Q�c�uχ�� ��t�f�x�:|���acces�? �+�=�O�a�s߅ߗ�Щ߻�������ne�ct to Network���%� 7�I�[�m�����(����ȘA��Ϻ���ϊ�!��`Int�roduction��t����������� ����(�OL^ p������� $5�_�P�*����VEditor5����
//�./@/R/d/v/5 T�ouch Pan�el � (re�commen�P) �/�/�/�/�/?#?5? G?Y?k?}?�̬P�^ �?�B�?OO/OAO SOeOwO�O�O�O�O�O <�O__+_=_O_a_�s_�_�_�_�_�_�Y�0�?�:�?o�?Eo Woio{o�o�o�o�o�o �o�o�OASe w������� ��+��_�_op�2o ������͏ߏ��� '�9�K�]�o�.���� ��ɟ۟����#�5� G�Y�k�}�<���`�¯ �������1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ��ώ��ϲ� �֯;�M�_�q߃ߕ� �߹���������%� �I�[�m����� ���������!���B� �f�(�*��������� ����/ASe w6������ +=Oas2� �V�����// '/9/K/]/o/�/�/�/ �/�/��/�/?#?5? G?Y?k?}?�?�?�?�? ����?O�COUO gOyO�O�O�O�O�O�O �O	__�/?_Q_c_u_ �_�_�_�_�_�_�_o o�? O�?Dono0O�o �o�o�o�o�o% 7I[m,_��� �����!�3�E� W�i�(o:oLo^o���o �����/�A�S�e� w���������~��� ��+�=�O�a�s��� ������ͯ������� ԏ9�K�]�o������� ��ɿۿ����П5� G�Y�k�}Ϗϡϳ��� ��������ޯ�� d�&��ߝ߯������� ��	��-�?�Q�c�"� t����������� �)�;�M�_�q�0ߒ� T߶�x�����% 7I[m��� �����!3E Wi{������ ���/��//A/S/e/ w/�/�/�/�/�/�/�/ ??�=?O?a?s?�? �?�?�?�?�?�?OO �6O�ZO/O�O�O �O�O�O�O�O_#_5_ G_Y_k_*?�_�_�_�_ �_�_�_oo1oCoUo go&O�oJO�o�o�_�o �o	-?Qcu ����|_��� �)�;�M�_�q����� ����xo�o�o���o 7�I�[�m�������� ǟٟ�����3�E� W�i�{�������ïկ ����ʏ��8�b� $���������ѿ��� ��+�=�O�a� ��� �ϩϻ��������� '�9�K�]��.�@�R� ��v��������#�5� G�Y�k�}����r� ��������1�C�U� g�y����������ߒ� ����-?Qcu ������� ��);M_q�� �����//�� ����X//�/�/�/ �/�/�/�/?!?3?E? W?h?�?�?�?�?�? �?�?OO/OAOSOeO $/�OH/�Ol/�O�O�O __+_=_O_a_s_�_ �_�_�_�O�_�_oo 'o9oKo]ooo�o�o�o �ovO�o�O�o�O#5 GYk}���� �����_1�C�U� g�y���������ӏ� ��	��o*��oN�� ��������ϟ��� �)�;�M�_������ ����˯ݯ���%� 7�I�[��|�>����� v�ٿ����!�3�E� W�i�{ύϟϱ�p��� ������/�A�S�e� w߉ߛ߭�l������� �ƿ+�=�O�a�s�� ������������� '�9�K�]�o������� ��������������� ,V�}���� ���1CU �y������ �	//-/?/Q/" 4F�/j�/�/�/? ?)?;?M?_?q?�?�? �?f�?�?�?OO%O 7OIO[OmOO�O�O�O t/�/�/�O�/!_3_E_ W_i_{_�_�_�_�_�_ �_�_�?o/oAoSoeo wo�o�o�o�o�o�o�o �O�O�OL_s� �������� '�9�K�
o\������� ��ɏۏ����#�5� G�Y�z�<��`ş ן�����1�C�U� g�y���������ӯ� ��	��-�?�Q�c�u� ������j�̿��𿲟 �)�;�M�_�qσϕ� �Ϲ����������%� 7�I�[�m�ߑߣߵ� �������߼���B� ��{�������� ������/�A�S�� w��������������� +=O�p2� ��j���� '9K]o��� d�����/#/5/ G/Y/k/}/�/�/`� ��/�/�?1?C?U? g?y?�?�?�?�?�?�? �?�O-O?OQOcOuO �O�O�O�O�O�O�O�/ �/�/ _J_?q_�_�_ �_�_�_�_�_oo%o 7oIoOmoo�o�o�o �o�o�o�o!3E __(_:_�^_�� ����/�A�S�e� w�����Zo��я��� ��+�=�O�a�s��� ����hz�� '�9�K�]�o������� ��ɯۯ���#�5� G�Y�k�}�������ſ ׿�����̟ޟ@�� g�yϋϝϯ������� ��	��-�?���P�u� �ߙ߽߫�������� �)�;�M��n�0ϒ� TϹ���������%� 7�I�[�m�������� ��������!3E Wi{��^���� ���/ASe w������� ��/+/=/O/a/s/�/ �/�/�/�/�/�/�? �6?��/o?�?�?�? �?�?�?�?�?O#O5O GO/kO}O�O�O�O�O �O�O�O__1_C_? d_&?�_�_^O�_�_�_ �_	oo-o?oQocouo �o�oXO�o�o�o�o );M_q�� T_�_x_���_�%� 7�I�[�m�������� Ǐُ돪o�!�3�E� W�i�{�������ß՟ 矦���>� �e� w���������ѯ��� ��+�=���a�s��� ������Ϳ߿��� '�9���
��.���R� �����������#�5� G�Y�k�}ߏ�N����� ��������1�C�U� g�y���\�nπ��� ��	��-�?�Q�c�u� �������������� );M_q�� ����������� 4��[m��� ����/!/3/�� D/i/{/�/�/�/�/�/ �/�/??/?A? b? $�?H�?�?�?�?�? OO+O=OOOaOsO�O �O�?�O�O�O�O__ '_9_K_]_o_�_�_R? �_v?�_�?�_o#o5o GoYoko}o�o�o�o�o �o�o�O1CU gy������ �_��_*��_�c�u� ��������Ϗ��� �)�;��o_�q����� ����˟ݟ���%� 7��X��|���R��� ǯٯ����!�3�E� W�i�{���L���ÿտ �����/�A�S�e� wω�H���l����Ϣ� ��+�=�O�a�s߅� �ߩ߻����ߞ��� '�9�K�]�o���� ��������Ͼ��2� ��Y�k�}��������� ������1��U gy������ �	-�����"� �F������/ /)/;/M/_/q/�/B �/�/�/�/�/??%? 7?I?[?m??�?Pb t�?��?O!O3OEO WOiO{O�O�O�O�O�O �/�O__/_A_S_e_ w_�_�_�_�_�_�_�? �?�?(o�?Ooaoso�o �o�o�o�o�o�o '�O8]o��� ������#�5� �_V�oz�<o����ŏ ׏�����1�C�U� g�y���������ӟ� ��	��-�?�Q�c�u� ��F���j�̯���� �)�;�M�_�q����� ����˿ݿ����%� 7�I�[�m�ϑϣϵ� ���Ϙ��ϼ����� W�i�{ߍߟ߱����� ������/��S�e� w����������� ��+���L��p��� F���������� '9K]o�@� �����#5 GYk}<���`�� ����//1/C/U/ g/y/�/�/�/�/�/� �/	??-???Q?c?u? �?�?�?�?�?��� �?&O�MO_OqO�O�O �O�O�O�O�O__%_ �/I_[_m__�_�_�_ �_�_�_�_o!o�?�? OOxo:O�o�o�o�o �o�o/ASe w6_������ ��+�=�O�a�s��� DoVohoʏ�o��� '�9�K�]�o������� ��ɟ�����#�5� G�Y�k�}�������ů ׯ�������ޏC�U� g�y���������ӿ� ��	��ڟ,�Q�c�u� �ϙϫϽ�������� �)��J��n�0��� �߹���������%� 7�I�[�m��ߣ�� ���������!�3�E� W�i�{�:ߜ�^����� ����/ASe w�������� +=Oas� ���������/ ���K/]/o/�/�/�/ �/�/�/�/�/?#?� G?Y?k?}?�?�?�?�? �?�?�?OO�@O/ dOvO:?�O�O�O�O�O �O	__-_?_Q_c_u_ 4?�_�_�_�_�_�_o o)o;oMo_oqo0OzO TO�o�o�O�o% 7I[m��� ��_���!�3�E� W�i�{�������Ï�o �o�o����oA�S�e� w���������џ��� ���=�O�a�s��� ������ͯ߯��� ԏ���
�l�.����� ��ɿۿ����#�5� G�Y�k�*��ϡϳ��� ��������1�C�U� g�y�8�J�\��߀��� ��	��-�?�Q�c�u� �����|������ �)�;�M�_�q����� �������ߜ߮��� 7I[m��� ������ E Wi{����� ��//��>/ b/ $�/�/�/�/�/�/�/ ??+?=?O?a?s?�/ �?�?�?�?�?�?OO 'O9OKO]OoO./�OR/ �Ov/�O�O�O_#_5_ G_Y_k_}_�_�_�_�_ �?�_�_oo1oCoUo goyo�o�o�o�o�O�o �O�O�o?Qcu �������� ��_;�M�_�q����� ����ˏݏ����o 4��oX�j�.������� ǟٟ����!�3�E� W�i�(�������ïկ �����/�A�S�e� $�n�H�����~���� ��+�=�O�a�sυ� �ϩϻ�z������� '�9�K�]�o߁ߓߥ� ��v��������п5� G�Y�k�}������ ���������1�C�U� g�y������������� ��	��������`"� ������� );M_��� �����//%/ 7/I/[/m/,>P�/ t�/�/�/?!?3?E? W?i?{?�?�?�?p�? �?�?OO/OAOSOeO wO�O�O�O�O~/�/�/ _�/+_=_O_a_s_�_ �_�_�_�_�_�_o�? o9oKo]ooo�o�o�o �o�o�o�o�o�O2 �OV_}���� �����1�C�U� g�x��������ӏ� ��	��-�?�Q�c�" ��F��jϟ��� �)�;�M�_�q����� ����x�ݯ���%� 7�I�[�m�������� t�ֿ��������3�E� W�i�{ύϟϱ����� �����ʯ/�A�S�e� w߉ߛ߭߿������� �ƿ(��L�^�"߅� ������������ '�9�K�]�߁����� ����������#5 GY�b�<��r� ���1CU gy���n��� �	//-/?/Q/c/u/ �/�/�/j���/? �)?;?M?_?q?�?�? �?�?�?�?�?O�%O 7OIO[OmOO�O�O�O �O�O�O�O�/�/�/�/ T_?{_�_�_�_�_�_ �_�_oo/oAoSoO wo�o�o�o�o�o�o�o +=Oa _2_ D_�h_����� '�9�K�]�o������� doɏۏ����#�5� G�Y�k�}�������r ������1�C�U� g�y���������ӯ� �����-�?�Q�c�u� ��������Ͽ��� ğ&��J��qσϕ� �Ϲ���������%� 7�I�[�l�ߑߣߵ� ���������!�3�E� W��x�:Ϝ�^����� ������/�A�S�e� w�������l������� +=Oas� ��h������� '9K]o��� �������#/5/ G/Y/k/}/�/�/�/�/ �/�/�/�?�@?R? /y?�?�?�?�?�?�? �?	OO-O?OQO/uO �O�O�O�O�O�O�O_ _)_;_M_?V?0?z_ �_f?�_�_�_oo%o 7oIo[omoo�o�obO �o�o�o�o!3E Wi{��^_�_�_ ���_�/�A�S�e� w���������я��� �o�+�=�O�a�s��� ������͟ߟ�� ��H�
�o������� ��ɯۯ����#�5� G��k�}�������ſ ׿�����1�C�U� �&�8���\������� ��	��-�?�Q�c�u� �ߙ�X���������� �)�;�M�_�q��� ��f�xϊ�����%� 7�I�[�m�������� ����������!3E Wi{����� ������> �e w������� //+/=/O/`s/�/ �/�/�/�/�/�/?? '?9?K?
l?.�?R �?�?�?�?�?O#O5O GOYOkO}O�O�O`/�O �O�O�O__1_C_U_ g_y_�_�_\?�_�?�_ �?�_o-o?oQocouo �o�o�o�o�o�o�o�O );M_q�� ������_��_ 4�F�
m�������� Ǐُ����!�3�E� i�{�������ß՟ �����/�A� �J� $�n���Z���ѯ��� ��+�=�O�a�s��� ��V���Ϳ߿��� '�9�K�]�oρϓ�R� ��v����Ϭ��#�5� G�Y�k�}ߏߡ߳��� ���ߨ���1�C�U� g�y���������� �϶�����<���c�u� �������������� );��_q�� �����% 7I��,��P�� ����/!/3/E/ W/i/{/�/L�/�/�/ �/�/??/?A?S?e? w?�?�?Zl~�?� OO+O=OOOaOsO�O �O�O�O�O�O�/�O_ '_9_K_]_o_�_�_�_ �_�_�_�_�?o�?2o �?Yoko}o�o�o�o�o �o�o�o1CTo gy������ �	��-�?��_`�"o ��Fo����Ϗ��� �)�;�M�_�q����� T��˟ݟ���%� 7�I�[�m����P��� t�֯�����!�3�E� W�i�{�������ÿտ 翦���/�A�S�e� wωϛϭϿ����Ϣ� �Ư(�:���a�s߅� �ߩ߻��������� '�9���]�o���� �����������#�5� ��>��b���N߳��� ������1CU gy�J���� �	-?Qcu �F���j�����/ /)/;/M/_/q/�/�/ �/�/�/�/�??%? 7?I?[?m??�?�?�? �?�?����0O� WOiO{O�O�O�O�O�O �O�O__/_�/S_e_ w_�_�_�_�_�_�_�_ oo+o=o�?O O�o DO�o�o�o�o�o '9K]o�@_� ������#�5� G�Y�k�}���No`oro�ԏ��$FMR2_GRP 1`���� �C4  B��p	 �p�0���F@ F�E���Q�F���C��L�F�Z!D�`�D��� BT��@����^�?�  x�����6������5�Zf5�ESΑ^�A�  ���BH��\���@�33@��� ����@�Q��@��g�]�Q����<��z�<�ڔ=7��<�
;;�*�<��^�8�ۧ�9k'V8���8���7ג	8(��~� ����=�(�a�L�����w�_CFG a�T0���ӿ������NO ��
F0+� 0���R�M_CHKTYP  �p	������ROMF�_MI�NL��s��x���7�X�SSB��b��� ���ϙu�����ϝ�T�P_DEF_OW�  �t	���I�RCOMK����$�GENOVRD_�DOm��q*�TH�Rm� dG�d0�_�ENB� 0�RWAVC��c���� �>�����v����^����.� �V��OU��i�3�q.��.�<u������,�z����sC�  D����l��2$�@��B�/��p1�m��ϑ�SMT���j��������$HoOSTC��1k�Κ���� M5C�t����v  27.0 =1��  e��B Tfx�
0�������	ano?nymous4 FXj|�r���������)
// ./@/R/�v/�/�/�/ �i/�/??*?<? N?����?�/�?� �?�?OO�/�?JO\O nO�O�?�O�/�O�O�O �O_S?�Ow?�?j_�O �?�_�_�_�_�_+Oo o0oBoTow_�O�O�o �o�o�o�o'_9_K_]_ _o5�_t���� �_����(�K}o �op����������o 13�$�gH�Z�l� ~������Ɵ؟��� �Q��D�V�h�z��� Ϗ�󏥯���;�� .�@�R�d��������� ����%���*�<� N�`ϣ���ǯ��ۿ�� �����&�i�J�\� n߀ߒߵ�7�����������"�o���ENT� 1l���  sP!��s�  u�a��������� 
������?�d�'��� K���o����������� *��Nr5�Y k�����8 �1n]�U�y ����/4/�X/ /|/?/�/c/�/�/�/��/�/?�/B?:QUICC0O?+?=?�?a41�?{?�?�?a4�2�?�?�?>O!ROUTER?OO-O��O!PCJOG��OjO!192�.168.0.1�0h?]3CAMPRYT�O�O!�E1�@_�FRTXO
__}_�C�NAME !~P�!ROBO�O��_S_CFG 1�kP� ��Auto-st�arted��FTP��a�Ϧ�Ao ��eowo�o�o�oF��o �o�o*o�oOa s���r��_oo �'Io�<�N�`�r� 5������̏ޏ��� �&�8�J�\�n�g�y� �ϝ�鏿�����"� 4�F�	�j�|������� ՟W������0�B� �������������ҿ �����ݯ>�P�b� tφϩ�+ϼ������� ��Y�k�}�/ߑς� ſ�߸������߱�� $�6�H�k�l��ߐ�� ��������-�?�Q�2� e�V���z�������s� ������
?���; dv������� %�9[�<N`r �G����� �&/8/J/\/n/�/� �����//?"? 4?F?X?/|?�?�?�? �?�/i?�?OO0OBO�TO�Z_ERR �m�Z\OlFPDUS_IZ  �0^0���D>�EWRD� ?�U�!� � guest�6�O�O __$_6_��TSCD_GRO�UP 3n�\ ��Q�9IFT|^$�PA|^OMP|^� |^_SH|^E�D�_ $C|^CO�Mn@TTP_AU�TH 1o{K �<!iPendCanBWMn�[�2�q�!KAREL:q*MoVohmKC}o��o�ou`VISI?ON SETfP�o�o�v!,rcP >hb�������~dCTRL �p{M6��1
1FFF9E3���$FRS:DE�FAULT[��FANUC We�b Server [�I��"d�O�D�я������+�jDWR�_CONFIG �qkU�Bc�[�lAIDL_CP�U_PCz��1B��� �� BH��M�IN��sQ��GNR_IOuA�B�0�H���NPT_SIM_�DOӖݛSTA�L_SCRNӖ ��ޚTPMODN�TOL�ݛ��RT�Y������` `EN�B�sS��OLN/K 1r{KxP�����ɯۯ������M/ASTEҐy�5����SLAVE �s{KH D��SRAMCACHE/�|A�"aO_CFGq������UO�`����CMT_OPz�ՒJ�ǳYCLp���t�_?ASG 1t`��A
 �6�H�Z�l� ~ϐϢϴ���������p� ��	�NUM�C5I
��IPn���RTRY_CNҿ���_UP_��A�����E ������u.)�  06��م��RCA_ACC �2vk[  R��� �) ��� 4@� 6���016��2?� ��#���  z�D���BUF�001 2wk[=� Bu��u0�Q��b��q�䂪�䑖䢖䱖�ª��і�����U����"��1�����Wu0*�J�@ku0H_W�z����������u0�\�@����u0"� S�u0#ߠQ����n�0u0Ch1ȫAn�Pn�an�p*n�n��n��n�M��f�پ��of`������,u0�rx�D��(gdu�0Pm��u0&@N��N�_�\p�����������Zx  Z�xR���R�&��&�&�&�&����S������s�2�����������t� x�������� ����������� ���������^�s��$�u�� ,��4��=��E���M�t� �T�t� �\�Ye��l�� t�q}�Y��y��q ��q��q��q��qx��qM��^����'�M���u0Z�����BH2����1�C8��3HA����	" 	"  	" $��,1" 5 1"= 1"E 1"M 1"�U ��\�e s=(lph�t��s�3����"�� �"�� ����"��� �"����"���2�� 2�2�2%� 2-�� 5�C2E�S 2U�� ]�2e�=�m� JPu�=���JP�� =���=���=�_4 ��=�� �� ���2 ���2���2���2���2 #�2##�Q$3# 2B5C#2BES#2BU c#�"e� 4t�&��;2xk[ 46�A�
�Q�P<J��D�AՒ���HIS}�zk[� �� 202?1-04-2J��S���� 9  +�>_P_b_t_�_�_�_��_�[L[SQ18-02-27_��_ok@��; Đ�B�b;c!�DQocopuo�o�o�[ZB��Xa6�_�o�o#o :���s.@Rdv.�ZY���X5�o���������B  7 �p�� 8 �:�9 ��2d��Ko�ZTI��X�"�������6��I��@: ��������(�:�LS���W19��n�����$����h�A6`pBd1B�pF�Ea�:d9�Db�q�S���XPK&Q���oI�[�m�9�9bF`K&Cc������ʯܯ�@�M� �O_;��7+P[�c�u��������� Ͽ��_�_?�)�;�)h��d9`�AdA`Y�I` Y�DχϙϫϽϫo�o ���)hqdp5�  �S�e�w߉ߛ߉� ��������+�=�+�*��c9�8'P_A�Y�
I�83�^Q�a�D�k� }�������ŏp��� 1�C�U�C�U������ ������a�ѐY� 5� �Y��a�9�Y���y� 2 �2���z�z�Y� ����������@�� �&�`%PT �������/@/�]J/\/%lB��iC7!f�DjC Ei/ �/�/�/�/�/��9/&?8?%l1bpAE?t?�? �?�?�?�߼�?OO (O:OLO^O'��19�	#�1f� I�1bQ�1b��O����O�O�O�� _4_F_X_j_|_j��|��_�_�_�_�_Ö �Qѐb��b�b  b9�b��bJo\oJ \�o�o�o��a�� �b�o�o&8&�I_CFG 2{�: H
Cy�cle Time~�aBusyDw�Idlzr�t�min={�q�Upvv|qRea}d�wDow�xܟۂqsCo�unt|q	Num� qr�s�={��`��q�PROGWr-|:D�0�u����������Ϗ�y �S�DT_ISOLCW  :�r�?�J23_DSP_�EN~ �>#�INC }��e��A   ?�=�?��<#�
�j�:�o u�������a��ȟ�OBK�C�,�FeU��G_GROUP 1~��< �� �j�Cy.�П?Dxd�m��`Q������̯@�����&�Dw���ڙG_IN_AU�TOdQ�#�POS�RE���KANJ?I_MASK��t��KARELMONG :(��by� ��(�:�L�@~²O�%�V�X��nŉ�ޛ�CL_Ld�NU�M0�����EYL?OGGING`?�j�U�F�LANGUAGE :�
��DEF�AULT �(L�GXq�V��r�~d�  8�p� ��`'�G  ��`�ۏ�;���
��(UT1:\\Ϧ� �ߵ��� �������!�8�E�W���(��#LN_DISP �M��x������OCTOL���aDz@��f���GBOOK �)ݹz�qz�z� Xr�k�}������������5Ӱs����	 -�t�*��/ُ`�+��_BUFF 2�^� A2�u v�ꂒ�w��� ��#,YPb ���������/��ZDCS �V�Y�n���#Dx^u��/�/�/�/6$IO ;2�B+ cp�/cp@���/??*?>? N?`?r?�?�?�?�?�? �?�?OO&O8OJO^O�nO�O�O�O�%ER_ITM��dD��O_ #_5_G_Y_k_}_�_�_ �_�_�_�_�_oo1o�CoUogo	��BSEVt�����FTYP����O�o�o�ovm��R�ST��4%SCRN�_FL 2��-@��g/gy�����TP�����b}�NGNAM,��`�
�2$UPS��G�Ip��U�B�_�LOAD�G �% �%DROP���MAXUALcRM�®� �U�9
��H�_PRM���� !���C����7������P �2�7� �q�	 �ol�W���{���Ɵ�� �՟���D�/�h� S�������¯���ɯ ۯ��@�+�d�v�Y� ������������߿� �<�N�1�r�]ϖ�y� ���Ϸ������&�	� J�5�n�Q�cߤߏ��� ��������"��F�)� ;�|�g�������� �������T�?�x� c����������������DBGDEF ��[!��_LDXDISA-��{�#MEMO_AP'��E ? �
 $x(�����������FRQ_�CFG ��6(A x'@�E��<[$d%m$�:������*�/� **:�����_�� ��+/"/4/a/X/j/ �/����/�@�/�/�/�/�',(�/>?�$,? i?P?�?t?�?�?�?�? �?OOOAO(OeOwO�^O�O��ISC 1� �� ����O�� )�O��2__V_�O�B�_MSTR ���myUSCD 1�o�N_�_J_�_�_o �_4oo1ojoUo�oyo �o�o�o�o�o�o0 T?xc��� ������>�)� N�t�_����������� ˏ���:�%�^�I� ��m�������ܟǟ � �$��H�3�l�W�i� ����Ư���կ��� �D�/�h�S���w���؛�Կj_MK'���]Y�$MLTA[RM&�-� 3" P�X� �METPUK ǲ����YNDSP_ADCOLr�& }�oCMNT�� ���FN���τ�FST�LI���ǁP ���^'�G�Y?�IԆ�P�OSCF����PgRPM��Y�ST���1��[ 4Q#�
��ϱ�����׿� ������7��+�m�O� a��������������E�/��SIN�G_CHK  ���$MODA%��K���DEV� 	N
	MC}:��HSIZEK�ǰ��TASK �%N
%$123456789  �2}�TRIG 1��[ l^`9n�=YP���5��~�EM_I�NF 1���`)AT&FVg0E0�+)�E0V1&A3&�B1&D2&S0�&C1S0=)�ATZ+fH@��:��bA�@/�'//K/]/  �/5GYk�/� ? 7/$?6?�Z??~?�? w?�?g/y/�?�/�/�/ 2O=?�/hO�?�OGOQ? �O}O�O�O
__�?@_ �?OO)O�_MO�_�O �_�_�Oo�_<oNo5o ro%_7_�o[_m__�o �_&]oJo� ;�����o��o �o�o�oX�|���� ��e֏�����0����NITOR�G� ?��   	?EXEC1˳s�U2y�3y�4y�5y�TC {�7y�8y�9˳t��rޔx�ޔ��ޔ ��ޔ��ޔ��ޔ��ޔ@��ޔ̒ޔؒޓ2�U2�2��2	�2�U2!�2-�29�2E�U2Q�3�3�3����R_GRP_S�V 1�  (�7񿩕�?����0B��r;�T�ǯo@�S&��
_Dς��9��ION_DB��|��Ǳ  ��e�����~��q��싷�  ��Ŧ�&�N   ������� h� }G��-ud1�����υ�PL_N�AME !�<��!Defa�ult Pers�onality �(from FD�)����RR2�� �1�L6�L�A�<��� d :҉ϛϭϿ������� ��+�=�O�a�s߅� �ߩ߻���������2��.�@�R�d�v�� �������<��� ��0�B�T�f�x���@�������޲���"��
���PJ \n������ ��"4FX' 9������� //0/B/T/f/x/�/ �/k}�/�/�/?? ,?>?P?b?t?�?�?�?�?�?�?�> H��6 H�b H�\���  �O1M�dC@PObM FO�O�G@�=�|C�Op�M�O�O C �H __ _2_P_V_t_�_��f��_�\��E	�`_�_o o�Q:�oA`�@oRodovn A�  �i �O�o�Lޱ�o�k�O �o'9$]H�J��R�� 1�4ɴ���R@ � �&�<��p @D� M �q?��s�q?���q�A��6Ez�  �q���;�	�l�r	 ��@� c0�ް!� ��p�� � � ��F��J��K� ��J˷�J�� �J�4�JR�<g|v�f0O����@�S�@�;�fA6A���A1UA���X{����=�N���f������T;f��X���ڀ��*  ���  �5Ó�>��p�H��?���?���#=�����ԏur`�f��q{��g���f���i�V���_(  ������Ȗt柉�	'�� � �I� �  ��eއ�:�È(�È�=���@����� <!�� �� �  ��qz���r��o�o����ү  �'覵��@!��p@�a�@��@���@��C�CR"��"��B�pC%�����@�r�������~n�������m;a;n�`@����D�u՟ҿ��������Q�c�E�UŔ�� �:�W  x�x?�ff�O�Ϙ�*�C �P���ˍ�8��<���>��x��q����0�P:�U�7�0�<0���>���|����<2�!<"7��<L��<`N�<D��<��,0h��ߴ��s��s Ҿ�`?fff?��?y&�аT@T����?�`?Uȩ?X�ᒩL��� �t,��t8��wW���� �ό�w�����������.��R���!�F��A���=���)����M����HmN �H[���G� F��HZE~ i�������  �oAK����� ���)���/�� %/7/�j/U/�/y/�/��/��M��"�i��C@�/?�/5? =8��??�F??j?��ç�s¬�-M�BH"��.���?,�[2�Y0X1�1@�Iܔ=@n��@��@: �@l��?٧]��? ��%��n�߱���=�=D��0O�B@��@�o�A�&{C/� �@�UXO�+J�8��
H��>���=3H���_�O F�6��G��E�A5�F�ĮE����O�@��fG���E��+E���EX��O�@>�\�G�ZE��M�F�lD�
�p�O�?E_0_i_T_ �_x_�_�_�_�_�_o �_/ooSo>owobo�o �o�o�o�o�o�o =(:s^��� ����� �9�$� ]�H���l�������ۏ Ə���#��G�2�W� }�h�����ş���ԟ ���
�C�.�g�R��� v��������Я	��� -��Q�<�u�`�r���zfB(hA4����h���൘�3���п��!4 �{x����!�0+#(Ϝ:��jbT�f�1?E�䴛|�Ђ� ���Ϯ��������i%P��P:�IVc߀��oߙ߄߽ߨف�� ��������9�$��"$<�N��r�����@v�H���&��e,��6�l�Z�|�����n)��������8�F
  2 H��6�&H�{�g\�b�&B�!�!� B��0
�0A� @�/��$�3@����l^�pUgy���$J0� � ��� 9T�%
 �� //+/=/O/a/s/�/��/�/�/�/�/^J� ���$����4��$MR_CABL�E 2�$� S� V�TP���@n�?�0F1�?0�)�0z Bz C[0n�OM�`B�����R6>n�:n�FG���n�??Q6 � B�� TO
��vr0��&��zn�n�E��O|�h�?�8� �� C� ]9h4��r0����.�~n��29�y��?�?�*\0�d� [@CW@j27��(�1n�=xP� 2I�/T3�OR˰O�O�O �O�O_�O�O"__*_ �_�_`_�_�_�_�_�_or5 +��_Qoco�uol�?o�o�o�ol��*�o** 3O�M �%9���zn�\�%%� 2345678'901%7u "R�Fqn�[@ �n��n�
Lw�nnot sent �j�zsW,�TE�STFECSALKGRI�gkʝd�td��q
�tG �P�n��"��'�9�K�� 9UD1:\�maintena�nces.xml�S���  ���DEFAULT�2GRP 2�	z  p�Sn��  �%1st� mechani�cal chec�kL}n��6��>�G�H�$r����������n��controller��7��Ic�8�J�0\�n���ϑM���n�"8��n�ȡϯH'�����*�<����Cٟn�����Y�����ҿ����ϒC��ge�. batteryς�W�H	���ϖϨϺ����ϑSupply? greasK���È�
�<���Hs�H�Z�l�~ߐ�zϑ �cabl��߾�g�
7���0� B�T��ؑ+�����Q�����������`�A$��@�hoo� �� ����������+� O� a�s�)Zl~�� ���'9 2 DV���{� ���
//k@/R/ �v/��/�/�/�/�/ 1/?U/g/<?�/`?r? �?�?�?�/�??-?O Q?&O8OJO\OnO�?�O �?�?�OO�O�O_"_ 4_�OX_�O�O�_�O�_ �_�_�_�_I_om__ To�_xo�o�o�o�oo �o3oEoWo>Pb t��o��o� ��(�:���p�� _����ʏ܏� �O� $�6���Z���~����� ��Ɵ��9�K� �o� D�V�h�z���۟���� ��5�
��.�@�R� ��v�ůׯ����п� ����g�<ϋ���r� ���ϨϺ�����-�� Q�c�8߇�\�n߀ߒ� �������)�;���"� 4�F�X�j�ߎ����� ���������m��� T���C���������� ��3�i�>��b t������/ S(:L^p��	 T~��� ��//&/8/J/\/ n/�/�/�/�/�/�/�/ �/?"?4?F?X?j?|? �?�?�?�?�?�?�?O�O0OBOTOfOxO � �?�  @� ��O�O�O���O__(_�*H_** ���@ zO|_�_�_b_�_�_�_�_��!__�_ Ko]ooo1o�o�o�oo o%o�o#5oA k}��o�oQ�� �E�1�C�U��� �a�����ӏ����	���e�w��
�$MR�_HIST 2���v�� 
 \��$ 2345678901����P�
BR��9������ ���?�Q�c��,��� ����t���ԯ��ί ;��_�q�(���L��� ˿��￦��%�ܿI�  �m��6ϣ�Z����������[�SKCFM�AP  �Uy��B�������ONREL  ��v�.�6��EXCFENB`�q
,��y�FNC���r�JOGOVLI�M`�dv����KE�Y`�����_P�AN_������RU�N����SFSP�DTYP��k��S�IGN`�r�T1M�OT��o��_C�E_GRP 1��.�~���O�� �÷���a������C� U��y�0�����f��� ����	��-?&c ����t�� ��Mq(��QZ_EDIT�]�(�Q�TCOM_�CFG 1�$������� 
�_/ARC_}�`���T_MN_MOD�E]���UAP�_CPL/��NO�CHECK ?^$� �� �/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?I��NO_WAIT_�L\���NT�ѭ$�3���1_E�RR��2�$�6ф �OEOWOiO�L<юO�O��53 OC�#M| ��,f���Bvſ����X�²�/C~���<�� ?���_�O?�7N�BPARAMB�.$���Df�_pb8ѫ_�[ = �� �_�_�S�_o(oo4o�^opoLo�o�o�kb���o�l}_n#UM_RSPACE!���b�GQt�$OD�RDSP#_��O�FFSET_CAqR�_/�vDIS��sS_A3 ARK�]�OPEN_FILE�p_���cq�PTION_IO������M_PRGw %3z%$*A�lS��sWO�p����C쀄���ꂗ  ;�?֞��g��	 ��Ȟ�����4�dpRG_DSBL  n��.�J��sRIE�NTTO_���Cٴ>�-�A �rUT�_SIM_D��+ҋBdpVhpLCT ��=���O}��=d\�_PEX; �n��RAT;' d������pUP �m��pw���� �|>�L��$PAL�2���>`�_POS_CCH�p��`�ZP2����L6�LA�W����oѯ �����+�=�O�a� s���������Ϳ߿� ��'�9ϵ�2��h� zόϞϰ��������� 
��CW�4�F�X�j�|� �ߠ߲���������*�wS$�4�5�4�Z�
BP G����������� ��&�8�J�\�n��� ��a�s��������� "4FXj|�� �������0 BTfx���� ���///_��g�Y/k-���c���/ �+�/�/�'>->-�o?�/3?�'tP(7R?H? Z?l?�?�?�?�?&0w�0�?L�D(4	`<?6OxHOZOA:�o<��xO�O�O�O�`A�  �I!?�O�__�] ?>_)_b_M___�_�_м_u����O�1����� ���$B@ ��؄��P @D� M a?�c�Q?<��a<�D�  Ezx0c�:�;�	l&b�	 �@�� 0�PP_` �
`� � � ��b��PH0#H���G�9G����G�	{Gkf����GΈK/�o�l�PC��1��`[�D	�? D@ D7g�n��d���  �O5��>(p`�4��(: B4�Bp{�!<�O��O��"���r'a�sW�Ao�R�ҧpߐ�p( W ��p�����_$��E	'� �� B�I� ��  ��E�F=����f�x���� <_`� �� � ��ف��8� b�__�GN=�� � 'N�(��aOpCR�`��`[pB`Cc�5�G� ���@�~�i���m?����G�MuAuN�@@<��*b7e ����4��X�C���𡃃���<�� :��a�tx?�faf�/į֯h� @���O�8<�3�A�>�׶q"a�J�pn��Px���uancnd؃>癙����u<2��!<"7�<L���<`N<D��<��,�o���c� c^��@?f7ff?�?& ��D�@T�2�?��`?Uȩ?X�B�:銒�'d�Ie v�g���Zd���ϵ� �������6�!�Z�l� Wߐߢ�y��߱���a���υ���D���HmN� H[�ArG� F��M���� ����������(�� %�^� _���K��� ��+���g�*<N �cu������Β���I={�C�O�s^?Ƀ�}���?yå�'c�'sqH�`�"xp��������:!@I�>}@�n�@��@:� @l��?���]/ ���%�n�߱����=�=D���n/� ��@��oA�&{C/�� @�U�/ ��+J8��
�H��>��=3�H��_�/ �F�6�G���E�A5F�Į�E���/� ���fG��E���+E��EX��?� >\�G��ZE�M�F�lD�
`8?/ �?n?�?�?�?�?�?�? O�?OIO4OmOXO�O |O�O�O�O�O�O_�O 3__W_B_{_f_x_�_ �_�_�_�_�_oo-o So>owobo�o�o�o�o �o�o�o=(a L�p����� ��'��K�6�H��� l�����ɏ���؏�� #��G�2�k�V���z��������韤"(�!4g�ퟦ����֕3�ϩ� ��!�4 �{:�L��!��0+#f�x�Z�j�b����1E���|��������"�P�F�4���P޲Px�����������׿¿��湿����A�,�Q�w�bϝ"$zό��� ������ߴ���@�.�d�R�ej�tߪߘߺ�������)����.���R�@�v��  2� H�6�&H�,����\��&B#�#B�  A� @ '�����"�4�F�W���߁���������T���$�� � �q�� ��%
 ��3EWi{� ������ܜ* ��b�����4�$PARA�M_MENU ?���� � DEF�PULSE�+	�WAITTMOU�T�RCV� �SHELL_�WRK.$CUR�_STYL��OPT���PT�B��C�R_DECSN�i�<,6/ H/Z/�/~/�/�/�/�/ �/�/?? ?2?[?V�SSREL_ID�  �����j5U�SE_PROG �%e%W?�?k3C�CR�|2��m�7_HOST !e#!�4O�:T���?�-C�?A/CiO�;_�TIME�|6�5~VGDEBUGz0�ek3GINP_F�LMSK�O�ITR\�O�GPGA�@ �L�p� [CH�O�HTWYPEbn�V? P?�_�_�_�_�_�_�_ oo?o:oLo^o�o�o �o�o�o�o�o�o $6_Zl~�� ������7��EWORD ?	e
 	RS�@^�PNS���s�JO!�TE<P@}�COL�3����3WL�0 ����	���5d�ATRA�CECTL 1�v��o v�U V������&����DT Q����S��D � t`�	 f��$Pf� f���f�v U����	��
d�Qu�ᦒc�uj�ur�Euz�u��	��������c�vj�vr�v
z�v��t��a�s��� ������͟ߟ��� '�9�K�]�o�������E��|0��U����U����E��! ����䡃2  ��,�>�P�����Ư د���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾�������� �*�<�N�`�r��������\� Ť� ����������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�U ���_ oo$o6oHoZo lo~o�o�o�o�o�o�o �o 2DVhz �������
� �.�@�R�d�v����� ����Џ����*� <�N�`�r��������� ̟ޟ���&�8�J� \�n���������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� ��_0�B�T�f�xϊ� �Ϯ����������� ,�>�P�b�t߆ߘߪ� ����������(�:� L�^�p������� ���� ��$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/�</N/X!�$PGT�RACELEN � W!  ���V �l&_�UP ���e��!� �!� �l!_CFG ���%�#V!� ���${#�/�(�- � ��%�"DEF�SPD ��,lU!~ �l IN� ?TRL ��-�!�8�%C1PE_CO�NFI� ��%'��!�$�)l WLID�#��-	�9�LLB 1�~7� ��$?B�  B4�3�& �5JOE�/ << T!?�1KPO1OHOjO�O ~O�O�O�O�O_�O�O@_L_2_T_�_�ZB �_�_�_�_3O�_"oo�'oXo�9GRP 1���<W!@� � �[�V!A?�x�D P�D�V�C2�� o�V d,D�i�i�1�0���0Wo)O�1�n��(s
�kB+pRq2�.hR�V!>'?oY>a�����~� =N�=R��3��0�i� T���x����Տ���<���  Dz0�9�V 
 �a��q����� ����ߟʟ��'���$�]�H���l�����)�W!
V7.10_beta1�$ܠ�B(�A�\�)A�G��aޡ>w������ޡ�A����ff�ޢA�p��AaG��Q�Q@�(��`� ��K�]�o����#Apأ�r�0�� ��Ϳ߿ڢU!��}����v�$��H�2ϝ:K�NOW_M  ��%�&�4SV �^�9��5N� ����f�9�$�6�o�(�"�m�3Mvc���} ��	�"V ����T���Pܽ�ߞ��פ�@ 1ߠ���(�wP�1+MRvcĥ�T~�D��u����OADB�ANFWD�ϡ3S�Tva1 1ś)��4�5�����& ��� �Q�D�V�h��� ������������
 O.@�dv������2�����V G�<%�w`3!3E��4bt����5������A6//,/>/��7[/m//�/��8�/�/�/��/��MA���d�3�'OVLD  �;�ߊ���PARNUM  �븆?�?��SCHS9 a5
�7�1�9��
EUPD�?�5uTO�%_CMP_��V0�����'��lDER_wCHKzE����0�ҎFwO�KRSg���Npa_MO���H_�O~�%_RES_G���;
8��oi_\_�_ �_�_�_�_�_�_o�_ /o"oSoFo9?+U6\F_xo+Ua�o�o�o -S��o�o�o-S  27-SZ Rqv-S � ���-S 0��<�-RV 1����ᾱ�@`z$�BT?HR_INRg�X1����dc�MASS6p� Z��MNo����MON_QUEUE ������@��U�$Nq@U�AN��ۈ�END��_��EXE ��6@BE����OPTIO���[��PROGR�AM %Պ%��.��?�TASK�_IU4g�OCFG� �Տ�?ɟ��D�ATA����@(�2��k�}����� ��^�ׯ�����ʯ�C�U�g�y�,�INFO���I���5�ҿ �����,�>�P�b� tφϘϪϼ�������@��(�:ߕ����I�� di���@DIT� ���߬���W�ERFLA�V���RGADJ Ή�/A�  ��?�@�w����� ��W�/�?���z��@'<@�9���%?h�0��dm�C�2�%糲+	H�l7�U�2�u?G�A ��t$���*��/�� **:���@������5,�'�����1��1W�9�Q����/�A� o�e�w����������� ��]G=O� s����5�� '�K]�� �/�����y/ #/5/c/Y/k/�/�/�/ �/�/�/Q?�/?;?1? C?�?g?y?�?�?�?)O �?�?O	OO�O?OQO OuO�O_�O�O�O�O �Om__)_W_M___�_ �_�_�_�_�_Eo�_o /o%o7o�o[omo�o�o�oN�	�<��*c Nt����Q�M����PREF ��%�����
��I�ORITY��܆�>��MPDSP������C�U������OD�UCT�������OG��_TG���钍ڂ�HIBI�T_DOA���TO�ENT 1Ӊ�� (!AF_I�NEm� �+�!�tcp+�S�!�udB�{�!iccmj�qXY��ԉ����)� 0��ߟ����ٟ� ��	�F�-�j�Q�c��� ��į��������$B�T�*����%����V����>}5o
�f��/	���������~��AG�,  ��o�D�V�h�(z��պ��Z뿺�������ϻ�i�EN�HANCE �u�s�A��d�P�7Մ~���������PORT_NUMn�������_C?ARTREP�Ĝ>�SKSTAm��oSLGS��ě��G�T�UnothingX�5�G��Y��{��TEMP �ڑ�e��e�_�a_seiban ���������"�� F�1�j�U���y����� ��������0@ fQ�u���� ���,P;t _������� //:/%/^/I/[/�/�/�/q�VERSI�L����  d?isablej�m�SAVE ۑ��	2670H7K55�(�/E?!@�0G?Y?|�}? 	�8w�$�o�;�?��e�?O"O4OFOTJ�<|?�Ot��5_�� 1�ě20�@r�e�O�O��g�pURGE�B掘�WFP�p�����W�3T�ѯ�W�RUP_DELA�Y ���&UR_?HOT %!vz��?߳_DUR_NORMAL�X���_�_�WSEMI�_�_;o�q_QSKIP�C�|��Cx�/�o�/�o�o�o �m}�o's�o!3E iW���w� ����/��S�A� c�������s�я���� ��ߏ�O�=�s��� ��]�����˟���>SRBTIF4T��RCVTMOU������/�DCR��C�^i ���aB4��B�q�(B[k@ϟ�k?�5�* ��{�m���#����A�ߒ��� $���o�ۯ�o <2�!�<"7�<L���<`N<D��<��9��O֯?�Q�@�u���������Ͽ�����)�;�o�R�DIO_TYPE�  �M1�G�ED��T_CFG ���KbBHSE��Xa2�� ���ȸ�����.� �ү D�/�h�S��ϙ�(o�� �o��ӟ�����;�)� _�M��m�ߴ�9�{� �������%��5�7� I���������a��� ����!E3i�� ���a�]�� �A/e��� mG���/�+/ /O/qv/�/G/�/C/ �/�/�/�/�/'??K? m/r?�/S?�?�?�?�? �?�?O�?!OW?}?nO�;���INT 2���Y���_�G;� ��O�K�+��OX�f�0 _[3O6_'OF_ H_Z_�_~_�_�_�_�_ �_o�_2oo*ohoVo �ozo�o�o�o�o�o
 �o.@&dR�v ���������<�"�`�N���!�EFPOS1 1�d�?  x\O҉ ���O����+�ŏ׏ �r�]���1���U�ޟ y�۟���8�ӟ\��� ����-�?�y�گů�� ��"���F��C�|�� ��;�Ŀ_�������� �B�-�f�ϊ�%Ϯ� Iϫ����ߣ�,��� P�b����Iߪߕ��� i��ߍ����L��� p���/����e�w� �����6���Z���~� �{���O���s�����  2����ze� 9�]���� @�d���5G ���/�*/�N/ �K/�//�/C/�/g/ �/?�/�/�/J?5?n? 	?�?-?�?Q?�?�?�? O�?4O�?XOjOOO QO�O�O�OqO�O�O_ �O_T_�Ox__�_7_ �_�_m__�_oo>o �_bo�_�o!o�o�oUc��2 1崏^opo �o(LRop� /��e���� 6����/���{��� O�؏s�������2�͏ V��z����9�K�]� ��������@�۟d� ��a���5���Y��}� �����ů��`�K��� ���C�̿g�ɿϝ� &���J��n�	��-� g��ϳ��χ�߫�4� ��1�j�ߎ�)߲�M� ��q߃ߕ���0��T� ��x���7����m� ������>������� 7�������W���{� ��:��^��� �ASe� �$ �H�li�= �a��/��� /h/S/�/'/�/K/�/ o/�/
?�/.?�/R?�/ v??#?5?o?�?�?�? �?O�?<O�?9OrOO��O1O�OUO�O�o�d3 1��o�O�O�OU_ @_y_O�_8_�_\_�_ �_�_o�_?o�_co�_ o"o\o�o�o�o|o �o)�o&_�o� �B�fx��%� �I��m����,��� Ǐb�돆����3�Ώ ���,���x���L�՟ p�������/�ʟS�� w����6�H�Z����� ����=�دa���^� ��2���V�߿z�Ϟ� ��¿��]�Hρ�ϥ� @���d����Ϛ�#߾� G���k���*�d��� ���߄���1���.� g���&��J���n� �����-��Q���u� ���4�����j����� ��;������4� ��T�x�� 7�[��> Pb���!/�E/ �i//f/�/:/�/^/��/�/?�OT4 1�_�/�/?�?m?�? �/�?e?�?�?�?$O�? HO�?lOO�O+O=OOO �O�O�O_�O2_�OV_ �OS_�_'_�_K_�_o_ �_�_�_�_�_Ro=ovo o�o5o�oYo�o�o�o �o<�o`�o Y���y��&� �#�\�������?� ȏc�u�����"��F� �j����)���ğ_� 蟃����0�˟ݟ� )���u���I�үm��� ���,�ǯP��t�� ��3�E�W����ݿ� ��:�տ^���[ϔ�/� ��S���w� ߛϭϿ� ��Z�E�~�ߢ�=��� a����ߗ� ��D��� h���'�a������ ��
���.���+�d��� ��#���G���k�}��� ��*N��r� 1��g���x8?045 1�;? ��1����� �/�/Q/�u// �/4/�/X/j/|/�/? ?;?�/_?�/�??�? �?T?�?x?O�?%O�? �?�?OOjO�O>O�O bO�O�O�O!_�OE_�O i__�_(_:_L_�_�_ �_o�_/o�_So�_Po �o$o�oHo�olo�o�o �o�o�oO:s� 2�V����� 9��]��
��V��� ��ۏv�����#��� � Y��}����<�ş`� r������
�C�ޟg� ���&�����\�寀� 	���-�ȯگ�&��� r���F�Ͽj�󿎿� )�ĿM��q�ϕ�0� B�Tώ�����߮�7� ��[���Xߑ�,ߵ�P� ��t��ߘߪ߼���W� B�{���:���^��� ������A���e�K]6 1�h�$� ^����� �$��H ��E~�=�a �����D/h �'�K��� 
/�./�R/��/ K/�/�/�/k/�/�/? �/?N?�/r??�?1? �?U?g?y?�?O�?8O �?\O�?�OO}O�OQO �OuO�O�O"_�O�O�O _|_g_�_;_�___�_ �_�_o�_Bo�_foo �o%o7oIo�o�o�o �o,�oP�oM�! �E�i���� �L�7�p����/��� S�������6�я Z�����S�����؟ s����� ����V�� z����9�¯]�o��� ����@�ۯd����� #�����Y��}�ϡ� *�ſ׿�#τ�oϨ� C���g��ϋ���&��πJ���n�	ߒ�x���7 1��?�Qߋ�	� ��-�3�Q���u��r� ��F���j������� �����q�\���0��� T���x�����7�� [��,>x� ���!�E�B {�:�^�� ���A/,/e/ /�/ $/�/H/�/�/~/?�/ +?�/O?�/�/?H?�? �?�?h?�?�?O�?O KO�?oO
O�O.O�ORO dOvO�O_�O5_�OY_ �O}__z_�_N_�_r_ �_�_o�_�_�_oyo do�o8o�o\o�o�o�o �o?�oc�o�" 4F�����)� �M��J������B� ˏf�������I� 4�m����,���P��� 럆����3�ΟW�� ��P�����կp��� ������S��w�����6����߷�8 1���l�~���6�!�Z� `�~�Ϣ�=ϟ���s� �ϗ� ߻�D������ =ߞ߉���]��߁�
� ���@���d��߈�#� ��G�Y�k�����*� ��N���r��o���C� ��g����������� nY�-�Q� u��4�X� |);u��� �/�B/�?/x// �/7/�/[/�//�/�/ �/>?)?b?�/�?!?�? E?�?�?{?O�?(O�? LO�?�?OEO�O�O�O eO�O�O_�O_H_�O l__�_+_�_O_a_s_ �_o�_2o�_Vo�_zo owo�oKo�ooo�o�o �o�o�ova� 5�Y�}��� <��`�����1�C� }�ޏɏ���&���J� �G������?�ȟc���ҿ�MASK +1���0�>�~�XNO  ��=�C�MOTE  �_�  ��_CFOG 휭��PL_RANG�������٦OWER� �����S�M_DRYPRG7 %��%��I���TART ��	�W�UME_PR�O&�8����_EX�EC_ENB  �����GSPD،�ΰָ�TD�B��RM��I_AIRPUR�� ��m�p��MT�_�T�����OB�OT_ISOLC�]��l�̥ȥ��N�AME ������OB_ORD_NUM ?	��i�H755  ��@�R�d���PC_TIME�OUT� x�S7232��1�`��� LTEA�CH PENDAaN�б�С��������Main�tenance /Cons�������"�ߒ�No Use�����@�R�d�pv�����NPOf�\��С����oCH_L������	���!U�D1:1���R�VGAIL!ц��������SPACE1 {2�`�
��@ХЩ�巓ΦТ�|m���< ���?�Y�Y���Kl C�|��������� %<�QrY `�d������Y )/@/�U/v/]/ �/������// 7/-?�/Q?r?�?k?�/ �/�/�/�/�??3?)O JO	O_O�OgO�O�?�? �?�?�?OOAO7__ [_|_�_e_�O�O�O�O �O�__=_3oToou_ �oqo�o�_�_�_�_�o o)o/Moe�] o�o�o�o�o�% G=�^����{��� ������!�S�9� ���o���g������2��� ��ݏ� ���%�W�Z���:�������Ưǟ3ڟ��� �"�ԯF�x�{���[� ��ҿ����4��� �1�C���g������@|��������	�5� .�@�R�d�߈ϺϽ߀ߝ������)�*�6 =�O�a�s߅�7���� ��$���5��J�K�7^�p����X��� ����E���5V-kl�8���������y �� f VwN���G ��� �ń
� �  �//1/ C/U/g/y/���-� ��/m�/ȁd0� /2?D?V?h?z?�?�? �/�/�.�:�?�;O? ?�?ZOlO~O�O�O�O �?�?�?�?O_5_(O :O�Oz_�_�_�_�_�_��O�O�O _"_4o `� @Ȁme�/ {oW__Y�a�UDo�o �o�_�j�o�o1Ca I��gq�� �����Q�c��� 7�i�����������Տ��ُ�\
�ol��A���*SYSTE�M*�V9.10�185 ��12/�11/2019 �A �� ��r��ӓSR_T  � � $ĐEN�B_TYP  � $RUNN�ER_AXS� �$HAND_LN�GTH�`�TH�ICK��FLIP�ґ�`$INTF?ERENCE��IF_CH��I�֑$�9�INDX�D�ĐG1POS   W�N�`��ANG`�x�_J�F��PRM`� �	�RV_DAT�AƑ  $���ETIME  ���$VALU�����GRP_ �  ��A  2 �SCő�	� �$I�TP_�� $7NUMڠOUِ	��TOT�
�DSP~!�JOGLIM� �$FINE_P7CNT@�CO���$MAX�TA�SK@�KEPT_�MIR=�]�PREsMTq�}�APLD���_EX�������t�@��PG��BRKHOLD�!��I_�  ڲ@��~�P_MADE��w�BSOC�MO�TN�DUMMY�163�SV_C�ODE_OPM�S�FSPD_OVR5D��R�LDL�O��ORZ�TPӐLEb[�F!�[�:�OV=�CSF��ᐓ�T�F�ƼA�a�UFRA��T�OOL@�LCHD�LYW�RECOVK��:�WSs�:��F=�ROM��I�_ᐮڐ @��S��N�VERT�OFSr;�CǠD�FWDt�x��p��ENAB���7�TR��`���E�_FDO��MB_�CM���B-�BLC_Mi�]��Ҫ�2S��VSTAA�$U�P�����G�׸�A�M����а��%� �_M��A�AM�A�1�OT$CA0�,�D�7�HBK���L�IO?�[�IQ�$PPAO�{�`���s��s�1�DVC_DB��F����쑼��A���1��%���3���+�ATIO� �h�K�U��/�/�P�ABF�T֒E�G�����E�:�_AUX~�SUBCPU�G�SIN_7Ў����P�1������FLA|��ݑHW_C1���j�����$AT�R���$UNIT������ATTR�I���G�CYCL�C�NECA!�F�LTR_2_FI�R�TARTUP_�CN`Ӷ�SIGN�O�LPS�2�1�_S�CTz�F_��F_��t��FSF����CHA��[���O��RSD/���/�P���s�_T��PRO8�|�p�EMP�=�"�T���ܐ����'DIAG�RAOILAC��p�M�LO��'�4�P�S-�@� i�+�%�P�R��SB�  z�C�� 	$ӯFUNC���RINS_TB���=��o�RA��`��7��a�E��WAR|q�8�BLCUR��$A+	((DA`��G(#%LD=� ?�h�o#��to#�TI��%�ܐ$�CE_RIA_S�WA�AF��P^�غ#��%T2\CK���CMOI���D�F_LE�_�PD��"LM��FA�H�RDYO��E�RG�t H� z���O 5MULSE� ���0�.�$JW�Jr����FAN_ALMsLV�Î1WRN�5�HARDאO�_O�,� �2�1STOd�Ƶ_���AU���R�(���_SBR ���5.�J���C_MPINFڐ��-De!8CREG@�N�V0l�$�۱DAL�_N��FL�����$M 2��7%�ܐ��8�ECM-�N0�YF�����G���SP�$R�$Y��Z�����ۡ��� ���EG!`
�?�F
QAR�0�'�20øU3 ��AXE$�R�OB!�RED!�W�R�߱_i]�SY�ܰDQᰋVS�WWRqI�V��STR �()��f�E��Ġ&T�o�1�B�P1��V5\c�OTOHAĠ�ARY�b]��ΡR�FI��h�$�LINK�!��3a�$EXT_�S1�r%U6�[aXYZ�2:ej7sfOFF9�2b)ZbNh`B����d�����cFI@ �g�A�7Ĩ9�_JL�¢d�?ch��0��T�[8�US��B�	qL2ArC7 ��DUtO�$V9pTUR�0!X�#zu!a(BX�P,�)wFL[`��@�P�p�|e�Y30�G� +1ĠKF�M�'Ł3��s�����a�ORQ.���x��s ��m�� �H��,�_AN]�OVEd���Mh  l��C~��C~��B}��0 {�B�|���{�~��h � ��e�u�����l�v��e�����C���.�E)RK��	tEЪ�$�E�A�ܐ�e�` gN!K�N!AX� ¢N!���4b��0�� Z1��o��`��r`��@�`��:p��qp��1�p ��:0��:0��:0Ǚ:0 י:0�:0��:0�:0��:0'�D�8�DEBU��$��3(�N�VbABNL�t�^�9VA�� 
��� �+���7�0�7�o7� a7�ra7��a7�:q7��qq�$Fp�"ۂ�cLA�B�b)�����GR�O: )r�<*�B_ ,��Tm��`�0��p*���1�AND�p�t�:�+�_e=��1Y�  *��A�Pm�!|�- ^`�NT�0ӟ�VEL�ل��L���SE�RVE���@ $��`�A]!��PO@ҹ ��`���@����!�@  ]$�TRQ�r
 �dtR
���"2��q I_ 	 l8���[ERR�bo�I,��لr�TOQلրLHP���R�� eG��%Ha��   ��REP  
 ,h��#�=�݁RA��? 2	 d��s��@��� �@�$r�� ����OC|?!�  d۟COUNT�Q��F�ZN_CFG	�# 4��aF3T���� ��ܣq ����AT��C/ �(�M��g2���Ճ{����FA� 䅻&��XdP��鐛��SQ��G�dQP~B���SHEL}@~Y� 5p�B_BAS��RS)R`F�^SS��!RM�1��M�2p�3p�U4p�5p�6p�7p�98��@�ROO�p���V ]`NL�ALsAB���FN�ACK�I%N�Tg �CU�0E0� 	_PUdq�2ZOU��P�aH-���� �P��TPFWD�_KARw�iAf�R�E��$0P/`U!w�QUE`I e�Up�r�0�1I�0�-�[`S��SF[aSEM3��A��0A��STYSO� 	�DI�}㸻���!_TMuCM�ANRQL[`EN�D�t$KEYSWITCH^s.��HEUpBEATmM�PEPLEv�(����UrF�s�S3DO_HOM�� O�1 EFA�PAR�a�vQ�P�EC��O01c���OV_Mxr� � IOCMGtd�A�	P,�HK�AG DXabG��U^�¹MP�W�WsFO�RCfCWAR 2���@.�OMP G @��c�0U�SEP3P1�&�@�$3�&Q4����O� L�"y��aHUNLO9 �\�4ED�1  ��SNPX_A�SZ� 0�@AD�D��$SIZ�fA$VA���M_ULTIP��.3�� A�! � �$H	/0��`BRS�}�ϱCrТ6FRI	Fu��S� �)��0{NFOODBU�P�~��5�3�9�ƽAfI�A�!$V�y�x�R�S|N��@ � L0Ə�TE�s8�:sSG%LZATAb�p&o�sCx᳍P[@STMT�q2�CPP�VBWe�\D�SHOW�Ev�BAN�@TP�`�wqs8���s8��r��V7�_Gv�� :p$PCD X�7���FB�!PX�SP� A U�AD�P��� �W�A00^�ZR� bW@� bW� bW� bW5`YU6`Y7`Y8`Y9`YA`YB`Y� bW��cV�@bWF`X7�$hlY(@�$h�Y@@$h�Y1�Y1��Y1�Y1�Y1�Y1��Y1�Y1i1i1�"i2_Y2lY2yY2��Y2�Y2�Y2�Y2��Y2�Y2�Y2�Y2��Y2�Y2i2i2B"i3_Y�p�xyY3�YU3�Y3�Y3�Y3�YU3�Y3�Y3�Y3�YU3�Y3i3i3"iU4_Y4lY4yY4�YU4�Y4�Y4�Y4�YU4�Y4�Y4�Y4�YU4�Y4i4i4"iU5_Y5lY5yY5�YU5�Y5�Y5�Y5�YU5�Y5�Y5�Y5�YU5�Y5i5i5"iU6_Y6lY6yY6�YU6�Y6�Y6�Y6�YU6�Y6�Y6�Y6�YU6�Y6i6i6"iU7_Y7lY7yY7�YU7�Y7�Y7�Y7�YU7�Y7�Y7�Y7�YU7�Y7i7i7"d���@P�U�# �߰e�
�A�2��� x #�R��@  ��M��RX9� ��Q_+�R��P��(�~ ��S/�C�D�^�_U�0i��"�YSL���� � L5Bj��4A7��D����&RVALU�j�% x1���F��IgD_L�3��HI���I�"$FILE_�L!�i$���S=A� h	�M�?E_BLCK�Z�|uAc�D_CPUsـM0s�A0u�$�6�-0Y�Z@FR  � PW-����0��LA�AS��������RUN_FLG ���� ���v�!���!���HF ��C���CA�T2x_LI�"�  ��G_O��� P_EDÍ"�@T2��c��k�9��nє0�0��B{C2LT �Q@` �(0�!c�FT�\��	TDC�A4�z���M�������T�H�0�!�#�$�Rx��0e ERVE�F�	F�5A�� ��  X -$q�LEN�~�	q��) RA� 2��W_�?���1q��2��MIOk�5S�0 I. �Z�����q���DE<�1LACE,":��CC3Z¶_MA�20>>TCVEfTXg
�|
@8RQ�QJ%AUM���J>JPR�}�2�`�@BP	0JKVK�A.)A.5A#�J�AF2JJ:JJBAAL2h:�hbAAf5#� NA1��XB G�L��a_�AA�ٱm�CF62�! `	�GROUP��vA�2$QN��C�3~�REQUIR1��0EBU�3m��$T 2 *!n�&8��50��" \� ��oAPPR  CLG��
$t�Ng(CLOD��w)S��)
��.u6# ���M �C 8� 2�$_MGA� �CLPN��(� R �'B{RK�)NOLD�&�@RTMOb�:
=�%Jb�4Pj  :�  B  �  �  6�W57W5hA���$�� "���Ax�7)A�3PATH�7��1�3�1���3� / #\�PSCA�� 7h"6�!INp�UC����Z0@C:PUM9HY��?�� @A��L�[J�0�[Jq0[@PAYLO�A7J2L�R_AN��CL�ЦI�A��I�A�%R_F2LgSHR@��ALO�D�~A�G=C�G=CACRL_��-E P)G�D�9H��G�$H�"NR�FLEXj#k�J��% PT"����E��W�A�kPp�& :}��� �W�T���0 ������F1�QEe Yg������(�bE2DVhz�� ��`x}t��m`@�x���QT�w^qXF���d�h% .�x1CUgkt�b������J�' �����	/����ATrf!� E�L�`��D�#(J/ &v* JE0CTR)A�maTN��@�'HA_ND_VBG�jQ����4( $�pF24�&���SW����TB�&)� $$M�@�)!��!�1 �#p��E2�A���@�&��<��-A�,���*A;A;G��+���*UD;D;P�0G�ІݩST�'�9�N8DY�e �&(�O� �@r��G�Q�G�A�G�t`�5P_5h5q5 z5�5�5�5�3 �R�4�* ��T�2 �a㵙!�ASYM$EeP F)K� L�A$O_B�X5@HD2=�4ĸ�ROdOvO�O�CJ��LR0�J�����Id_�VI��ؙ#!�V_UN���6�W��AJN�|�N��LR�U _ԃ�]� $YR03_E_$���[TcS α��3HR���+���L}P]"DI0#O#�������,) g�V�I9�AV1S P�s`^�^�v`��ϰ�`�� - � ɑME�a��y���`�T�PT��Հ�0����V ��������T��� $�DUMMY1q1o$PS_p`RF2`���$���PFL�A�YP���?$GLB_T��1���]!S��aq�}��. XT '�1ST��* SBR�0M�21_V&"T$S/V_ER�@O��w��CLK�w�A�`OlS� �GL�EW��/ 4���$Y
��Z��W���Aœ�Az�9BΥ0��U.��0 �pN����$GI��}$>�� /������1 L���}�$F��ENEA�R�`NwcFd	�`T�ANCwbͱJOG�&`H0 2Ӑ$JOINT�"���޽�MSET�3 E EJ�a�S������4� �n`U�a?�* LOCK_FO�@Б�oBGLVt�GLTEST_XMj N�EMP� &"2I�� $U�P��9`#20* ��X1#̐4� X/y�CE�&�y $KAR$qM>%�TPDRA����VEC`�� I�UX2]HE T�OOL9c�V8dR�E�IS3�U�6�z1m`ACH� / 3��O@����3g��% SIZ"  @�$RAIL_BO�XE���ROB�O)?���HOW�WARVQH!��!ROLM�n%ԁ$"p�6 a`�0O_F��!��HTML5D�)A��!�15�*5�R�O�R6�1`��� ґ��OU�7 d��T/`�J�$��� $PIP*N �p�6"!`X� �P?CORDED� 
@L� a XT*0) �� �O`� 8 D 0�OB|�N�� ��7v1��/�v2��P�S;YSv1ADRO� ���TCH� 9� ,�pEN	�QA
_�4݁0����VWVA|�: Ǥ ����PR�EV_RT��$�EDIT(FVSHWR�c�G@�b��%�D��O�^DW�?$HEAD����4x@��0CKE�����CPSPD�FJM%P�0L�ϰR�`;�;~0{Q�6I3SO�C��NE�P���OTICK9c��M�Q�Ͳ�CHNY�< �@�0�AᅗA_GP8&V-&�PSTY�2!LOK���B"R�P_= t 
#@G�5S%$A=c�SE�!$D�9`���M�r�P&�&VSQU�x,e��TERC�����אS�>   o���p��q�``1O����{`IZ����PR\0�Db��A0PU;�Te_DYOi�0XS� K�AXIs`�#]UR��cP�O P�6����_��2ET�bP��0	�Ԑ� 
�sPA,����9'[�) ��SR��?l�P�!���/u�Ay �/u*�/s8�/sH�uu j�uuz�uu���u�}����u�|���yC
��}C��}�ϕϧϹ�5�SS}C3� @ h��cDS4P/���SPJ�&��ATx� �UaP��B��ADDRESz�B3@SHIF�^O_2CHO��1�IR���TUR�I��� A�CUSSTO�d��V�I>�AB�2��8c�
2�
 BV1da~�C 	\a�8�rPC�a�P��C��b�bR�6������TXSCRE�Ex2D��QTICNA��# Ӕ�A8�a��ٰE T�A�� 8b�1��n� ��a�2�b�/@RROS�~ �0��@�o�� UE�DF# ���1
�S��1'RSMPwgUe0�P抡�S_��=� ����ȧ=õaC����� 2EΐUE�մGD���D`GM�T��Lp��a~�O��� BBL_ W���~�H �rPJ�O��V�LE�a�N ��`�RIGHj�B�RD��ہCKGR�����Tf0����WIDTH#T@�b)!�j�i�I� EY���}�I
2� m VR6 @aBACKTQ�Ś����FOS1�L[AB_q?(��I �$URT!E�"��ް��H@� J 	8��~ _wA�h�R���s(����U�)O�~�KP�����Uv���Ry!LUqM�ØfՀERV!1RR�Ph �L���`�GEI�O�`l2�@LIP��bE�Pf�)%�@v�3؆�3�  2�50�60�70�8��R��?`h ���� !�Sv�PKݱUSR��OM <a���U�(�FO�PR�I�am  ���TR�IP2!m�UN+DO;�N �P ��ye`!xeS�P�`�P �Oc���CaG �PT� T��^�OS��s�R�`F�J��Z�P��������6Th�P	U�Z�Q���ãҜ5UJ�OFF([�R�_���O)� 1�P���;�Q��GU�1P:�V�Q�`���SUB6R���SR	T��tSR}� #csOR ��RAU(p"��T���7��_&@�D�T |1p�8OWN|M��4$SRCQ��Ҡ�PD(&rMP�FIMTl��`ESP Pab����eA���p����A@
�U `���WO[p�4a�PC�OP��$�`O�_`- ��1�WA3@CF�� Z��"��@l"+� V�SHADOW�`��?_UNSCA���ʴDGD!�1E�GAC�8�K�V�CWp`
�W� �,"w1�S$NEAR�c�Q#+�C0^cDRIV6f�aC_V/P��@m D��?MY_UBY��k�yV��UR��P�eA�� "P_MT"mLZkBM]�$�@7DEY�3EX7�^��MU�@X]�V$��cUS���`�_R鑠����
�R���G�pP�ACIN�A�PRG �$�"�"��"ң��RE}�遚�c�8H�"@X �� �G�P��� @�IR��@Y��?�ӱ���	�qaREb#SW&� _A�!�`W#B`�O��ہA�^3/rE"��UeP�d��J+HKjRZ��v:�P0&q[0%��3EAP�7�� j�^5�IMRC]V
�[ ��OvPMj�C��	�2��#�2REF6�F�6�1 M0���c50���:FAJ FAKhE�6�?_ �:�H�;�pS��N'�ap����I�\ �GR��ӵ`�м�PO�U4W�"Vk )W 5U�2��$Ԑ��C`,�Y��U�2Q{��ՀULj�Z_ C�O~��[H EPNTZ�T��U���V���SQPL��U#�U����W���VIA_܃��] ��`HD<����$JO��6���$Z_UP)L�W�Z|pW!e�Q�PSp�0�_LI��$EPEQ��k�a�Q�Ǒ΁��΀G\m�^�� 0���aw� ޴�CACHLO :A�d�aI �i��� 1-CI`MI�FHa�eqT�p�f�K$HOj�z�`COMM���Ot�wWӲ�S&�T7 VP�"@�mrO_SIZwtZ� `rx!asw���MP�zWFAI!`G�4�`sAD�y�MRET�r|wGP��> & �ASYNBUF�VRTD�%�|q���OL�D_��A�W6��PC��TU7#�`yQ{0	�ECCU�(�VEM� �e���gVIRC�q9�!���%�_DELA�#&Q���AG5�RK!X#YZ̠��K!W1���8A��򱦀TN8"I�M߁8������eGRWABB��Yb" �e��_e��LAS���A�a_GE�e` u�&��;���T/S&N` ���%I���"ņ��BGf�V5��PaK� ǆ�aWGI��	N#�`2�A@��`�q�q�a+�aS�p�fN\:�]�LEX��b�@����;��Nq��I? ��-|�� |�.$�3Pk��- �"c��b��t�Ŀ��a�ORD�����Q��w�RN�d� $MPTIT�� �C��F�VSF����e  -�[�QfK UR�3]�SM!�sf+���ADJ��N%�PZD>�g DƨBaAL+`�p�Ab�PERIs`��MS7G_Q9�$}q�u���b��h+�"�g�xJ`�3p�XVR#��in�b�T_OVR~i���ZABC��aj�";�s/@
 i��Z]�#�k+�=$L��-B�ZMPCEF��lH���A��®�LNKc�
^�M�K!��m $x,q�0��CMCM� �C�C���DP_=A+A$J����Dbq���� �� `����
D�F�UX���UXE]!f��	� ]��]�oс�oё���FTFsQӾ�A9�b�n {�}�����YJ`D�� o�Y�R�pU�$H�EIGH�#"�?(�MP�.A����Dp� � EX�$B�QPx �SHIF,�s��RVI`F��/B|�0�C`�dTF @{"�������WuD��_TRACE��V�A�^� PHER� q ,MP�)�;��$R�!p�� ����F�W\� 6�S�>F��  S�x�(2p������s����r�����	��U�C��ADC��=l6�R  d�� �ZD �Qx0C�����l�l0�| �r6�V��@ 2F����� D� P �����	�	F�,: $ZH~l��� ���� //D/2/ h/V/x/�/�/�/�/�/ �/
?�/??.?d?R? �?v?�?�?�?�?�?O �?*OONO<OrO`O�O �O�O�O�O�O�O__ 8_&_H_n_\_�_�_�_ �_�_�_�_�_�_4o"o XoFo|ojo�o�o�o�o��o�oF��$SAF�_DO_PULS C�G��k�$qp����|k���5qR ��`�XP�B\�\�[������(�s��[� �� ������*�<�`N�`�r������  ��2��[�[�d�������rs�� @������*��܉�� � 6��/_ @J�TY J����������T D��������)� ;�M�_�q����������˯ݯ��~�����M�_�$��sNR�;��f����p���
�t��Di��q��  � ����R�q |ulq���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w������S��G����� ��0�B�T�f�x��� ��������������@"4FK��b0E� ҳD�ܽ����� �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?��?�?�? �?�?�?�?	OO-O�� QOcOuO�O�O�O�O�O �OLz��!_3_E_ W_i_{_�_�_�_�_�_ �_�Yoo,o>oPobo to�o�o�o�o�o�o�o (:L^p��������ø� �Ǔ�6�H�Z�l�~� ������Ə؏����  �2�D�V�d�#�m�\����������i�	12345�678ݲh!B�!ܺTz1!���
��.�@�R� d�v�������"�ïկ �����/�A�S�e� w���������ѿ��� ���)�;�M�_�qσ� �ϧϹ��������� %�7����m�ߑߣ� �����������!�3� E�W�i�{��L߱��� ��������/�A�S� e�w������������� ��+=Oas ������� '9��]o�� ������/#/ 5/G/Y/k/}/�/N�/ �/�/�/�/??1?C? U?g?y?�?�?�?�?�? �?�/	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_BS��]_�o_�?�_�_�_Ԛ�Cz  Bp�z �  ��2��� } �X
g_�  	��R2U_ <oNo`oro�l��\�+o�o�o�o�o" 4FXj|��� �������oB� T�f�x���������ҏ �����,�>�P�b� t����������Qa:�R<Ք ˕a?  ������#a#at  ��P#�;���`�$�SCR_GRP �1*P�3 � ��R� �U	 _����� �����Qԑ�U������pٯǯ ��]�`6��C�,����m���C����lLR �Mate 200�iD 56789�0!`LRM|� 	LR2D ��~�
1234���Ц�d��hbճ ���}�ݣ}��cԑ����ѡ�	j4�F��X�j�|τ���#H���Ē�}��πį������̦<��1���A���e��WV��Vh�`,R��  -��B��Pư߮���Ԫ�A�P��  @��0�ժ�@����� ?4���H�P'������F@ F�` Q�Y�P�}�h���� ���������ʩ������J�5�G�Y�k�B� y������������ =(aL�p���o�
'�����W�`�.4�@4�>'�}�4̧@��n�PȄ����ݣT_��A���ߒ���aĲ�1  
/1/C/Q*!f(r/$�/S/�P�#
b�/ �/�/� ?�/$?,4]��ECLVL���1�����>1L_D?EFAULTF4������0~Z3HOTSTRf=��z2MIPOWEKRFE0�Ur5�4oWFDOg6 r5�=2RVENT 1�M1M1�3 L!�DUM_EIP�,?H�j!AF�_INEf0+O3D!'FTOZN!O~O9!�ϣO �mO�O�!RPC_MAIN�O�H��O_�C'VIS�O�I�_b_o!TPUPPUY_�IdQ_�_!
PM�ON_PROXY�_Fe�_�_uR�_M�f�_Fo!RDMO_SRVGoIg5o��o!R���oHh,�o�o!
�@MoL�i�o*!RLSgYNC+Qy8>v!ROS O�|��4e�!
CE>wPMTCOM�F�k��!	�rCO�NS�Gl�Z�!}�rWASRCao�FmI���!�rUSB��Hn���O �Uc���?�d�+����O���s�П87RVI�CE_KL ?%��; (%SVCPRG1ן�	�2�$��3G�L��4o�t��5�����6��į�7���H��/�*�97�<�� �od������9��� �a�ܿ������� ,��ٯT���|�� )����Q���6�z��� 6����6�ʿD�6�� l�6�ϔ�6�Bϼ�6� j���6����6���4� 6���\�^�
�ܟ�� �������.������ 8�#�\�G���k����� ����������"F 1X|g���� ��	B-f Q�u����� /�,//P/;/t/�/ q/�/�/�/�/�/�/?�?(?L?7?p?�_D�EV �9��UT1:|?�0GRP 2
�5����bx 	� 
 ,�0x?�?�2 �?OO@O'O9OvO]O �O�O�O�O�O�O�O_ *__N_5_r_�_�?�_ __�_�_�_o�_&o8o o\oCo�ogoyo�o�o �o�o�o�o4�_) j!�u���� ����B�)�f�x� _�������������M �,��P�7�t�[�m� ����Ο�����(� �L�^�E���i����� �ܯ�� ����6�� Z�l�S���w������� �ѿ���2�D�+�h� ��]Ϟ�U��ϩ����� ����@�R�9�v�]� �߬ߓ��߷������� *��N�`�G��k�� ����������&�8� �\�C�����y����� ����C���4F- jQ������ ��B)fx _�������� /,//P/7/t/�/m/ �/�/�/�/�/?�/(?p?!?^?e3d �e6	L?�?�?�?�?�?�?�OK%�O5O<C���NA�1NE^OlG VO�OzO�O�O�O�I"O _JI�O4_"_X_F_h_ j_|_�_�O�__�_o �_0ooToBodo�_�_ �o�_�o�o�o�o, P�ow�o@�< �����(�jO� ����p�������܏ ʏ �B�'�f���Z�H� ~�l�������؟��� >�ȟ2� �V�D�z�h� ����ůׯ�������� .��R�@�v�����ܯ f�п������*�� Nϐ�uϴ�>Ϩϖ��� ��������&�h�Mߌ� ߀�nߤߒ��߶��� .�T�%�d���X�F�|� j��������*�� ���.�T�B�x�f��� ����������� *P>t�����d ����&L �s�<���� ��/T9/K//$/ �l/�/�/�/�/�/,/ ?P/�/D?2?T?V?h? �?�?�??�?(?�?O 
O@O.OPOROdO�O�? �O O�O�O�O__<_ *_L_�O�O�_�Or_�_ �_�_�_oo8oz__o �_(o�o$o�o�o�o�o �oRo7vo jX �|����*� N�B�0�f�T���x� ������&����� >�,�b�P���ȏ���� v���r�����:�(� ^�����ğN�����ȯ ʯܯ� �6�x�]��� &���~�����Ŀƿؿ �P�5�t���h�Vό� zϰϞ����<��L� ��@�.�d�R߈�v߬� ����ߜ����<� *�`�N���߫���t� ��������8�&�\� �����L��������� ����4v�[��$ �|�����< !3��T�x ����8�,/ /</>/P/�/t/�/� �//�/?�/(??8? :?L?�?�/�?�/r?�? �? O�?$OO4O�?�? �O�?ZO�O�O�O�O�O �O _bOG_�O_z__ �_�_�_�_�_�_:_o ^_�_Ro@ovodo�o�o �o�oo�o6o�o* N<r`���o� ���&��J�8� n������^���Z�ȏ ���"��F���m��� 6���������ğ��� �`�E����x�f��� ����������8��\� �P�>�t�b������� ��$���4�ο(��L� :�p�^ϔ�ֿ������ �π���$��H�6�l� �ϓ���\��ߴ����� �� ��D��k��4� ������������� ^�C����v�d����� ������$�	���� ��<r`����� � �$&8 n\������ �/� /"/4/j/� �/�Z/�/�/�/�/? �/?r/�/i?�/B?�? �?�?�?�?�?OJ?/O n?�?bO�?rO�O�O�O �O�O"O_FO�O:_(_ ^_L_n_�_�_�_�O�_ _�_o o6o$oZoHo jo�o�_�o�_�o�o�o �o2 V�o}� FhB���
�� .�pU�����v��� �����Џ�H�-�l� ��`�N���r������� ޟ ��D�Ο8�&�\� J���n�����ݯ� �����4�"�X�F�|� �����l�ֿh��� ��0��Tϖ�{Ϻ�D� �Ϝ����������,� n�Sߒ�߆�tߪߘ� �߼����F�+�j��� ^�L��p������ ��������$�Z�H� ~�l������������ �� VDz�� ���j���� 
R�y�B� �����/Z� Q/�*/�/r/�/�/�/ �/�/2/?V/�/J?�/ Z?�?n?�?�?�?
?�? .?�?"OOFO4OVO|O jO�O�?�OO�O�O�O __B_0_R_x_�O�_ �Oh_�_�_�_�_oo >o�_eowo.oPo*o�o �o�o�o�oXo=|o p^����� �0�T�H�6�l� Z�|�~���Ə��,� �� ��D�2�h�V�x� Ώ�ş������� 
�@�.�d�����ʟT� ��P�ί�����<� ~�c���,��������� ʿ�޿�V�;�z�� n�\ϒπ϶Ϥ����� .��R���F�4�j�X� ��|߲������ߢ��� ���B�0�f�T���� ����z���������� >�,�b������R��� ����������:|� a��*����� ��Bh9xl Z�~���� >�2/�B/h/V/�/ z/�/��//�/
?�/ .??>?d?R?�?�/�? �/x?�?�?O�?*OO :O`O�?�O�?PO�O�O �O�O_�O&_hOM___ _8__�_�_�_�_�_��_@_%od_nQ�$S�ERV_MAILW  nUd`�Jh�OUTPUTYh�oP@NdRoV 2�V  g`� (�Q4o�oNdS�AVEzlhiTOP�10 2�i d j_ 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ����U��eYP�oKcFZN_CFG �Ugc�d�a�eT�?GRP 2^��a� ,B   A���nQD;� B����  B4�c�RB21�fHELLW��U�f�`�ou���%RSR��)�b�M��� q�����ο��˿��@(��L�7�pρ��Ͽ�  �a%@�����Ϗ͓���oP1��������Ǫ��2oPd����ɦHKw 1׫ � �߃ߕߧ��������� ��%�7�`�[�m��������ìOMM� ׯ�ȢFT?OV_ENBYd�a��iHOW_REG�_UI7�LbIMI_OFWDL�����l�WAIT4� ��v���t`X��d��wTIMX������VAX`��l�_UNcIT3��iLCQ�WTRYX��eN`�MON_ALIA�S ?e��`heo�����
t ��#�GYk }�:����� �/1/C/U/g//�/ �/�/�/l/�/�/	?? -?�/Q?c?u?�?�?D? �?�?�?�?O�?)O;O MO_OqOO�O�O�O�O vO�O__%_7_�O[_ m__�_�_N_�_�_�_ �_o�_3oEoWoioo zo�o�o�o�o�o�o /A�oew�� �X������ =�O�a�s�������� ͏ߏ����'�9�K� ��o���������b�۟ ������"�G�Y�k� }�(�����ůׯ鯔� ��1�C�U� �y��� ������l����	�� ƿ?�Q�c�uχ�2ϫ� �������Ϟ��)�;� M�_�
߃ߕߧ߹�d� ������%���I�[� m���<�������� ���!�3�E�W�i�� ��������n����� /��Sew�����$SMON_�DEFPROG �&����� &*S?YSTEM*��� 	�RECA�LL ?}�	 �( �},cop�y frs:*.�dt virt:�\temp\=>�192.168.�1.15:630�0 F416 6��l~�}
xy�zrate 61 ,>P��/���0 ��b/�t/�/�tpdiosc 0+/0 =/�O/�/�/?�tpconn 0 �/��/�/_?q?�?� 11 ,?>?P?�?�?O��.!md:pick.tp��;�?�aOsO�ONdrop -O?OQO�O�O_/�O�0�?�Oa_s_�_�?1 )?=_O_�_�_o_)_ �_�_^opo�o�_�_9o Ko�o�o o%o�o�o l~�o�o5GY ��!���h� z����1�C�U���� 
��O�O��ӏd�v��� �>�?�Q������� ����ϟ`�r������� ;�M�ޯ���'��� ˯\�n�������7�I� ������#���ǿٿ j�|Ϗ���3�E�W��� ���ϱ�����f�x� �ߝ�/�A�S������ ߭߿���b�t��� ��=�O�������)� ����^�p������9� K����� �%����� l~����5GY ��!���h z��1CU�� 
/���d/v/�/ �-/?/Q/�/�/?/ +/�/�/`?r?�?�/�/@;?M?�?�?O�7!��frs:orde�rfil.dat~0�mpback;���0�?jO|O�!�b:*.*6O�>PO�O�O�_T�$SNPX�_ASG 2����,Q�� P 0 '�%R[1]@X�0_WY?��%W_ �_f_�_�_�_�_�_�_ o�_7oo,omoPowo �o�o�o�o�o�o�o 3W:L�p� ������ �'� S�6�w�Z�l������� �Ə����=� �G� s�V���z���͟��ן ��'�
��]�@�g� ��v��������Я�� #��G�*�<�}�`��� ����׿��̿��� C�&�g�J�\ϝπϧ� �϶�������-��7� c�F߇�j�|߽ߠ��� ��������M�0�W� ��f���������� ���7��,�m�P�w� �������������� 3W:L�p� ����� ' S6wZl��� ��/��=/ /G/ s/V/�/z/�/�/�/�/ ?�/'?
??]?@?g? �?v?�?�?�?�?�?�?�#ODTPARAM� ,U6Q ��	�'JP'Dj@'H~D�-P�POFT_KB_?CFG  C2U�SOPIN_SI/M  ,[sF�O��O�Ov@=@RVNO�RDY_DO  �}E�ERQST_P_DSB�NsB�U_aX=@SR ��I � &�@E�STa_�^�T�CT�OP_ON_ER�R_;B�QPTN ��E�P��C�RRING_P�RM�_0RVCNT?_GP 2�E�A�@x 	Q_Po@`>owobo�olWVD%`�RP 1LI�@ �axI�g�o�o�o EBTfx��� ������,�>� P�b�t�������яΏ �����(�:�L�^� p���������ʟܟ�  ��$�6�]�Z�l�~� ������Ưد���#�  �2�D�V�h�z����� ��¿����
��.� @�R�d�vψϯϬϾ� ��������*�<�N� u�r߄ߖߨߺ����� ����;�8�J�\�n� ������������ �"�4�F�X�j�|��� ������������ 0BTf���� ����,S�Pbt����bPRG_COUN�P�D��R�ENB�o�M��D/_U�PD 1{[T  
�BR/d/v/ �/�/�/�/�/�/�/? /?*?<?N?w?r?�?�? �?�?�?�?OOO&O OOJO\OnO�O�O�O�O �O�O�O�O'_"_4_F_ o_j_|_�_�_�_�_�_ �_�_ooGoBoTofo �o�o�o�o�o�o�o�o ,>gbt� �������� ?�:�L�^��������� Ϗʏ܏���$�6� _�Z�l�~�������Ɵ������_INF�O 1@%9& H�	 �c��N���r�@
U�@CIy=���t���Bv�ſ��X��n²�C~��⒭>�� @g�� A��`=��` >`� >����� C	����	(>B���hC3��9!�C2������@�D"(>�N���a�3��]��2���Y?SDEBUG�A ���d))Q�SP_�PASS�B?~c�LOG =�]J!  �����  �%!�UD1:\��#���_MPC��@%�#ϒ@!̱A� @!�SAV ���y�ظ�вC�׸SV��TEM_TIM�E 1��K � 0  $��$Q~C�%�C�+���MEMBK  @%%!����%�7�G��X|& � @G���iߎߞ�b�d������^� y�@����*�<�v�T��f�x������ � ������
��.�@�R�d�v��e�������� ����(:L^ p������� ��SK������@RdX�� "��2sߣ�`�  ���������%/7/I/8[/O�u$� �u/���ߴ/�/�/���/��?'?9?K?]?o?�� s?�?���?�4^�?�? �?OO/OAOSOeOwO �O�O�O�O�O�O�O_�_)�T1SVGU�NSPDy� '�c��4P2MODE_LIM ��dg�0T2=P]Q���/UASK_OPTGIONX��g��Qw_DIr�ENB���c��QBC2_GRP 2#c���_��� C�c(\BCCFG !�[�~���p!Ekem` eo���o�o�o�o�o�o �o?*cN` �������� �;�&�_�J���n�����ˏݏ�Ȍ��ɏ *�<����r�]����� ��H�ڟԯ����� ,��P�>�t�b����� ��ί������:� (�J�p�^��������� ܿʿ�� �6��� J�\�zόϞ���ϰ� �������.�@��d� R߈�v߬ߚ߼߾��� ���*��N�<�r�`� ������������ �$�&�8�n�\���H� ����������|�" 2XF|��n� ����0 fT�x���� �/�,//P/>/t/ b/�/�/�/�/�/�/�� 
??:?L?^?�/�?p? �?�?�?�?�? O�?$O OHO6OlOZO|O~O�O �O�O�O�O_�O2_ _ B_h_V_�_z_�_�_�_ �_�_�_�_.ooRo? jo|o�o�o�o<o�o�o �o<N`.� r������� &��J�8�n�\����� ��ȏ���ڏ���4� "�D�F�X���|���ho ʟܟ������B�0� R�x�f���������� ү���,��<�>�P� ��t�����ο���� �(��L�:�p�^ϔ� �ϤϦϸ������ȟ *�<�Z�l�~��Ϣߐ� ��������� ���D� 2�h�V��z���� ����
���.��R�@� b���v����������� ��N<r(� �����\��8&\Fz�$�TBCSG_GR�P 2"F��  �z 
 ?�  � �������5/�/Y/k+~�$�_d@ ��!?z	 HBLk(z�&~j$B$  C��0�/�(�/�/Cz�/(=�A�k(333?&�ff?��i%A���/m?80 k(�1͎6S5�0DHp?�=@�H0j%K1�5j$�1D"N!�?�?�?�?;O J�(I&�(nE�OLO^O �O�O�O�O�O_ [�H�:Q	V3.0�0�	lr2d S	*\PTTyk_f*_ �Q�I �Pt]�_  �_�_�[~J2�%�=Qo~�UCFG 'F�� �"j��Lb�ROlwl� wo�o�jO�o�o�o�o �o=(aL^ �������� �9�$�]�H���l��� ��ɏ��Ə���#�� G�Y��� d�v���2� ����˟�ܟ� �9� $�]�o�����N����� ۯƯ��zf6�B F�H�Z���~�����ؿ ƿ����2� �V�D� z�hϞόϮϰ����� ���
�@�.�d�R�t� �߈߾߬����ߴ� ���>�`�N��r�� ���������&��� 6�8�J���n������� ��������"24 F|j����� ��B0fT �x�����/ �,//P/>/`/�/0� �/�/�/l/�/�/?? ?L?:?p?^?�?�?�? �?�?�?�?O O"OHO ZOlO&O|O�O�O�O�O �O�O_�O_ _2_h_ V_�_z_�_�_�_�_�_ 
o�_.ooRo@ovodo �o�o�o�o�o�o�o *�/BT�� �������8� J�\��l��������� ڏ����ʏ4�"�X� F�h���|�����֟ğ ���
���T�B�x� f���������Я��� ��>�,�b�P�r�t� ����6Կ�����(� �8�^�Lς�pϦϔ� ������ ߾�$��H� 6�X�~ߐߢ�\�n��� ������ ��D�2�T� z�h���������� ����
�@�.�d�R��� v������������� *N`
�x�� F����$ J8n��Pb� ���/"/4/F/ / j/X/z/|/�/�/�/�/ �/?�/0??@?f?T? �?x?�?�?�?�?�?�? �?,OOPO>OtObO�O �O�O�O�O�Ol�_ ._�O_L_^_�_�_�_ �_�_�_ oo$o6o�_ ZoHojolo~o�o�o�o �o�o�o2 VD fhz����� ��
�,�R�@�v�d� ��������ΏЏ�� �<�*�`�N�����@_ ����ҟ|���&�� 6�8�J���n�����ȯ گ�����"��F�0��  l�p� �p���p��$TBJ�OP_GRP 2�(8�� _ ?�p�	��ڣ�*���@���@�� 0��  �� � � � �{p� @l����	 �BL  ~ �Cр D�����<��E�A�S�<��B$�����@��?�33C�*���8œϞ� ��2�T�����;�2��t��@���?���zӌ�-�A5�>�Ⱥ�� ������l�>�~�a�s�;��pA�?�f�f@&ff?�ff�ϵ�8� ��L����}������:v,����?L~�}ѡ�DH���5�;�M�@�33`�����>��|օ��8���`ự�	�D"��������`�r��|���"�9�� ����g�v��x��נ� ������������0 (V�b��`���p�C�p��	���	V3.�0�	lr2d��*b��k�p{� E8� E�J� E\� E�n@ E��E��� E�� E��� E�� E�h� E�H E�0 E� Eϒ��� E��� E�x E�X� F��D�  D�` E�_P E�$�U0�;�G�R��^p Ek�u�������(��� E�����X� 9�IR4! DH%�
z�`/r"p��v#Ѭ߱/��ESTPARSI d������HR� ABLEW 1+��J p���(�' �k)�'B�(�(o�w��'	�(E
�(�(5p��(��(�(K!�#RD	I�/��??(?:?L?^5�4O�?�;�?�?�O O2N�"S�?��  �:�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo���@�O ��7�isO�O�O�OU?�g?y?�?�?�8�"pbN�UM  8�*����x� J K ��"_CFG ,�Y{s�@��IMEBF_TT�!u��� �vVERI#�a�v��sR 1-�+' 8mp�k�� ;��o  ��� ,�>�P�b�t������� ��Ώ�����(�:� ��^�p���������ʟ ܟ� ��$�6�H�Z� l�~�������Ưد� ��� �2�{�V�h��� ������¿Կ���
Ϥ�"�q_Sq�v@�u�� MI_CHAN�w �u u�DBGLV���u�u�!x��ETHERAD �?�%���v ��������(x�RO�UT�p!WJ!�*�H��SNMAS�K���s��255.��N�ߖߨ�N� �OOLOFS_D�I� BŪ�ORQCTRL .�{>Cw/&�T�J�\�n� ������������� �"�4�F�X�j�z���������#PE_D�ETAI����PG�L_CONFIG� 4Yyiq���/cell/$C�ID$/grp1���;M_q�9C� ߮����� ,>Pbt�� ����/��:/ L/^/p/�/�/#/�/�/ �/�/ ??�/6?H?Z? l?~?�??1?�?�?�?�?O O�n}�?VOhO zO�O�O�Oq���O�M��?__1_C_U_g_ �?�_�_�_�_�_�_t_ 	oo-o?oQocouoo �o�o�o�o�o�o�o );M_q �� ������%�7� I�[�m�������Ǐ ُ�����!�3�E�W� i�{������ß՟� �����/�A�S�e�w� �������ѯ������ �User View )	�}}1234567890J�\�n����������5�	̿��0�2=���� �2�D� V�h�ǿٿ7�3�� ���������o�1�߾4��j�|ߎߠ߲���#���߾5Y��0�B�@T�f�x��ߙ�߾6� ��������,���M�߾7�������������?�߾8u�:L�^p������ �lCamera;�1�0BT2BE�~� �H�����//�  ���f/x/ �/�/�/�/g�/�/? S/,?>?P?b?t?�?�����?�?�?�?O O,O�/PObOtO�?�O �O�O�O�O�O�?�7X� �O>_P_b_t_�_�_?O �_�_�_+_oo(o:o Lo^o_�72+�_�o�o �o�o�o�_*<N �or�����so ���a�(�:�L�^� p��������܏�  ��$�6���7t�͏ ��������ʟܟ�� � �$�o�H�Z�l�~��� ��I��7(	9�� �� $�6�H��l�~���ۯ ��ƿؿ���ϵ�ǧ9��O�a�sυϗϩ� P������Ϙ��'�9ߠK�]�o߁�
	�0 ߼���������� :�L�^�߂���� ����ߕ�� ���5� G�Y�k�}���6���� ��"���1CU ���I+������ ����1C�g y����h�յ; X//1/C/U/g/ �/�/�/��/�/�/	? ?-?��![�/y?�? �?�?�?�?z/�?	OO f??OQOcOuO�O�O@? ��k0O�O�O	__-_ ?_�?c_u_�_�O�_�_ �_�_�_o�O��{�_ Qocouo�o�o�oR_�o �o�o>o);M_<qm  i� �������0�xB�T�f�   v ~������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ�j�  
`(  ��p( 	  ���B�0�f�Tϊ� xϚϜϮ��������t,���� ��o q߃ߕ��������� ��c`�=�O�a�� ���������&�� �'�n�K�]�o����� ����������4�# 5GYk������ ���1C �gy����� ��	/P-/?/Q/� u/�/�/�/�/�//(/ ??)?p/M?_?q?�? �?�?�/�?�?�?6?O %O7OIO[OmO�?�O�O �O�?�O�O�O_!_3_ zO�Oi_{_�_�O�_�_ �_�_�_oR_/oAoSo �_wo�o�o�o�o�oo �o`o=Oas ���o�o���8 �'�9�K�]�o���� �����ۏ����#� 5�|�Y�k�}�ď�����şן���B�"�@ A�*�<�N��$�����+frh:�\tpgl\ro�bots\lrm�200id��_m�ate_��.xml
���Ưد����` �2�D�V�F���`� ��������Ϳ߿�� �'�9�K�b�\ρϓ� �Ϸ����������#� 5�G�^�X�}ߏߡ߳� ����������1�C� Z�T�y�������� ����	��-�?�V�P� u��������������� );R�Lq� ������ %7NHm�� �����/!/3/tE.g��� $��r�<< p� ?�E+�/E/�/�/�/ �/�/?�/?<?"?4? V?�?j?�?�?�?�?�?��?�?
O8OF��$�TPGL_OUT?PUT 7P�P�_ h tE �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o�tEh �=@2345?678901Lo^o po�o�o�o�cF�Io�o �o�o/�o3e w���Ez}�� ���'���]�o� ��������O�ŏ��� �#�5�͏C�k�}��� ����K�]������ 1�C�۟Q�y������� ��Y�ϯ��	��-�?� ׯ�u���������Ͽ g�ݿ��)�;�M�� [σϕϧϹ���c�u� ��%�7�I�[���i� �ߣߵ�����q����@!�3�E�W���HA}c!�������������@�j/�.�p* ( 	 1oc�Q���u� ��������������) M;q_��� ����7%�GI[��?f� f &��-�#/5/ /Y/k/9j��/�/H/ �/�/�/�/?,?�/0? b?�/N?�?�?�?�?�? >?�?O�?OLO^O8O �O�O�?|O�O�OvO _ _�O_H_�O�O~_�_ *_�_�_�_�_�_ol_ 2oDo�_0ozoTofo�o �o o�o�o�o�o.@ dv�o^��X ����*���`� r����������ޏ<� N��&���2�\�6�H� �������ڟt�Ɵ� "���F�X���@���(� z�į֯�����j��� B�T��x���d����� �0���Ϣ��>�� *�tφ�俪ϼ�VϨ��������(�:��)�WGL1.XML���o��$TPOF?F_LIM ����}�Nw_SV��  �����P_MON �8������2y�STRTC�HK 9�������VTCOMP�AT��6��VWV_AR :��Y�.�� � q�������_DEFPROG %�ه%������ISPLAY���ޡ��INST_MSK�  �� ��I�NUSER,���L�CK5���QUIC�KMENY���SC�REx��7�tpsc��5��h���ҩ�_��ST*����RACE_CF�G ;��Y����	z�
?���HNL 2<��`� ��L^p������
��ITE�M 2=8 ��%$123456�78901  �=<)Oai  #!ow��3� z��A//w)/ ��v/��/��/�/ M/=/O/a/{/�/�/�/ U?{?�?�/�??'?9? �?]?	O/OAO�?MO�? �?�?qO�O#O�O�OYO _}O�OX_�Os_�O�_ �__�_1_�_og_'o �_7o]ooo�_{o�_	o o�o?o�o#�oG �o�o�oSk�� ;�_q:��U�� y�������%��I� 	�m��?�ŏ��Ǐُ ���w�!�͟��i� )�������+�՟���� ���ůA�S�e��7� ��[�m�ѯy����п +��O��!υ�7ϩ� ����߿��ϯ����� K���oρϓ�߷�c� �ߛ��Ͽ�#�5�G��� ��}�=�O��[����� �����1����g��P���f���S��>>k��  �k�� ����
 ���������UD�1:\&��}�R_GRP 1?�� 	 @ ��q�m��������  �&�J5nY?�   �������/ �//'/]/K/�/o/��/�/�/�/�/�/	�9�?%?{�SCB ;2@�� tq? �?�?�?�?�?�?�?O�q�UTORIAL� A��LOv�V�_CONFIG B����	�O[M�OUTPUT yC���@���O �O__1_C_U_g_y_ �_�_�_�_�_�A�O�_ oo1oCoUogoyo�o �o�o�o�o�_�o	 -?Qcu��� ���o���)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����+� =�O�a�sυϗϩϻ� �������'�9�K� ]�o߁ߓߥ߷����� �����#�5�G�Y�k� }����������O �E�O'�9�K�]�o��� ���������������� #5GYk}�� �����1 CUgy���� ���	/-/?/Q/ c/u/�/�/�/�/�/�/ �/?/)?;?M?_?q? �?�?�?�?�?�?�?O ?%O7OIO[OmOO�O �O�O�O�O�O�O_ O 3_E_W_i_{_�_�_�_ �_�_�_�_o_/oAo Soeowo�o�o�o�o�o �o�oo+=Oa s������� ��&9�K�]�o��� ������ɏۏ����>�����0�B� ,��m��������ǟ ٟ����!�3�E�W� i��������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sτ��� �ϻ���������'� 9�K�]�o߀ϓߥ߷� ���������#�5�G� Y�k�}�ߡ������ ������1�C�U�g� y�������������� 	-?Qcu�� ������ );M_q��� ����//%/7/ I/[/m//��/�/�/ �/�/�/?!?3?E?W?�i?{?�;�$TX_�SCREEN 1}DD�,���}ipnl/��0gen.htm��?�?�?OO%O���Panel soetup)L}�)O@jO|O�O�O�O�OXO NO�O__1_C_U_�O y_�O�_�_�_�_�_�_ n_�_-o?oQocouo�o �_,o"o�o�o�o )�oM�oq��� ��BT��%�7� I�[�� ������Ǐ ُ���t�!���E�W��i�{�������>UA�LRM_MSG k?�9��0 �� �*��5�(�Y�L�}� p�������ׯʯ�����ӕSEV  ��Q�ђECFoG F�5�1�  �%@�  }A��   Bȍ$
  ��#�5��ƿ ؿ���� �2�D�V��h�v�]�GRP 2�Gg� 0�&	 �����ӐI_BB�L_NOTE �Hg�T��#l�"�0�!s��¿DEFPROݐ%� (%�:ߖ  (�a�L߅�pߩߔ��� �������'��K����FKEYDATA� 1I�9��p 	v��&�ϰ����������,(�+��$��OINT  ]�3�5� OOK T���{�b�NDIRE�CT���� CHO�ICEN���F�UC�HUP����F�RE INFOO aH�l���� ��9 ]o� ��/fr�h/gui/wh�itehome.pngp�������  �point�*/</N/`/r/�//look"g /�/�/�/�/�/*indirec/�4?F?X?j?|?.clos�'?�?�?�?�?�O*touchup$?<ONO`OrO�O.arwrg#?�O�O �O�O_�H#_5_G_Y_ k_}_�__�_�_�_�_ �_o�_1oCoUogoyo �oo�o�o�o�o�o	 �o?Qcu�� (������� ;�M�_�q�������~ ��ӏ���	��-�4� Q�c�u�������:�ϟ ����)���;�_� q���������H�ݯ� ��%�7�Ư[�m�� ������D�ǿ���� !�3�E�Կi�{ύϟ� ����R�������/� A���S�w߉ߛ߭߿� ��`�����+�=�O� ��s�������\� ����'�9�K�]�������������v��������#5WiC,U�M���� ��<N5rY ������/� &//J/1/n/�/g/�/ �/�/�/���/?"?4? F?X?g�|?�?�?�?�? �?�?w?OO0OBOTO fO�?�O�O�O�O�O�O sO__,_>_P_b_t_ _�_�_�_�_�_�_�_ o(o:oLo^opo�_�o �o�o�o�o�o �o$ 6HZl~�� ����� �2�D� V�h�z������ԏ ���
���.�@�R�d� v��������П��� ���/<�N�`�r��� ������̯ޯ��� &���J�\�n������� 3�ȿڿ����"ϱ� F�X�j�|ώϠϲ�A� ��������0߿�T� f�xߊߜ߮�=����� ����,�>���b�t� �����K������ �(�:���^�p����� ������Y��� $ 6H��l~��� �U�� 2D�V-�X�-�������}���,�/
/�/./ /R/d/K/�/o/�/�/ �/�/�/??�/<?#? `?r?Y?�?}?�?�?�? �?�?O�?8OJO)�nO �O�O�O�O�O��O�O _"_4_F_X_�O|_�_ �_�_�_�_e_�_oo 0oBoTo�_xo�o�o�o �o�o�oso,> Pb�o����� �o��(�:�L�^� p��������ʏ܏� }��$�6�H�Z�l��� ������Ɵ؟�����  �2�D�V�h�z�	��� ��¯ԯ������.� @�R�d�v���_O���� п�����*�<�N� `�rτϖ�%Ϻ����� ���ߣ�8�J�\�n� �ߒ�!߶��������� �"��F�X�j�|�� ��/����������� ��B�T�f�x������� =�������,�� Pbt���9� ��(:�^ p����G��  //$/6/�Z/l/~/��/�/�/�/���+}�������/@?=�/7?I?#6,5O z?-O�?�?�?�?�?�? �?O.OORO9OvO�O oO�O�O�O�O�O_�O *__N_`_G_�_k_�_ �_���_�_oo&o8o G/\ono�o�o�o�o�o Wo�o�o"4F�o j|����S� ���0�B�T��x� ��������ҏa���� �,�>�P�ߏt����� ����Ο��o���(� :�L�^�ퟂ������� ʯܯk� ��$�6�H� Z�l���������ƿؿ �y�� �2�D�V�h� ���Ϟϰ��������� �_�.�@�R�d�v�}� �߬߾��������� *�<�N�`�r���� �����������&�8� J�\�n�����!����� ��������4FX j|����� ��BTfx ��+����/ /�>/P/b/t/�/�/ �/9/�/�/�/??(? �/L?^?p?�?�?�?5? �?�?�? OO$O6O��8K�����aOsO�M]O�O�O�F,�_�O�__�O2_ D_+_h_O_�_�_�_�_ �_�_�_�_oo@oRo 9ovo]o�o�o�o�o�o �o�o*	�N`r ����?���� �&�8��\�n����� ����E�ڏ����"� 4�ÏX�j�|������� ğS������0�B� џf�x���������O� �����,�>�P�߯ t���������ο]�� ��(�:�L�ۿpς� �Ϧϸ�����k� �� $�6�H�Z���~ߐߢ� ������g���� �2� D�V�h�?������ ������
��.�@�R� d�v������������ ����*<N`r ������ �&8J\n� �������"/ 4/F/X/j/|/�//�/ �/�/�/�/?�/0?B? T?f?x?�??�?�?�? �?�?OO�?>OPObO tO�O�O'O�O�O�O�O __�O:_L_^_p_�_h�_�_}��[�}�����_�_�]�_o)of,Zo ~oeo�o�o�o�o�o�o �o2VhO� s�����
�� .�@�'�d�K�����y� ��Џ����'_<� N�`�r�������7�̟ ޟ���&���J�\� n�������3�ȯگ� ���"�4�ïX�j�|� ������A�ֿ���� �0Ͽ�T�f�xϊϜ� ����O�������,� >���b�t߆ߘߪ߼� K�������(�:�L� ��p�������Y� �� ��$�6�H���l� ~���������������  2DV]�z� �����u
 .@Rd���� ���q//*/</ N/`/r//�/�/�/�/ �/�//?&?8?J?\? n?�/�?�?�?�?�?�? �?�?"O4OFOXOjO|O O�O�O�O�O�O�O�O _0_B_T_f_x_�__ �_�_�_�_�_o�_,o >oPoboto�oo�o�o@�o�o�o��{��������ASe}=��sv, ���}����$�� H�/�l�~�e�����Ə ؏����� �2��V� =�z�a�������ԟ�� ��
���.�@�R�d�v� ���o����Я���� ���<�N�`�r����� %���̿޿��ϣ� 8�J�\�nπϒϤ�3� ���������"߱�F� X�j�|ߎߠ�/����� ������0��T�f� x����=������� ��,���P�b�t��� ������K����� (:��^p��� �G�� $6 H�l~���� ���/ /2/D/V/ �z/�/�/�/�/�/c/ �/
??.?@?R?�/v? �?�?�?�?�?�?q?O O*O<ONO`O�?�O�O �O�O�O�OmO__&_ 8_J_\_n_�O�_�_�_ �_�_�_{_o"o4oFo Xojo�_�o�o�o�o�o �o�o�o0BTf x������ ��,�>�P�b�t����]���]�����ÏՍ����	��,��:��^�E� ����{�����ܟ�՟ ���6�H�/�l�S��� ����Ư���ѯ� � �D�+�h�z�Y���� ¿Կ�����.�@� R�d�vψ�ϬϾ��� ����ߕ�*�<�N�`� r߄�ߨߺ������� ���8�J�\�n�� ��!����������� ��4�F�X�j�|����� /����������� BTfx��+� ���,�P bt���9�� �//(/�L/^/p/ �/�/�/�/���/�/ ? ?$?6?=/Z?l?~?�? �?�?�?U?�?�?O O 2ODO�?hOzO�O�O�O �OQO�O�O
__._@_ R_�Ov_�_�_�_�_�_ __�_oo*o<oNo�_ ro�o�o�o�o�o�omo &8J\�o� �����i�� "�4�F�X�j������ ��ď֏�w���0� B�T�f������������ҟ���� ���>� ���!�3� E��g�y�S�,e��� ]�ί�����(�� L�^�E���i������� ܿÿ ����6��Z� A�~ϐ�wϴϛ����� �/� �2�D�V�h�w� �ߞ߰��������߇� �.�@�R�d�v��� �����������*� <�N�`�r�������� ��������&8J \n����� ���4FXj |������ /�0/B/T/f/x/�/ �/+/�/�/�/�/?? �/>?P?b?t?�?�?'? �?�?�?�?OO(O�� LO^OpO�O�O�O�?�O �O�O __$_6_�OZ_ l_~_�_�_�_C_�_�_ �_o o2o�_Vohozo �o�o�o�oQo�o�o
 .@�odv�� ��M����*� <�N��r��������� ̏[�����&�8�J� ُn���������ȟڟ i����"�4�F�X�� |�������į֯e������0�B�T�f��$�UI_INUSE�R  ������� � g�k�_MENHIST 1J���  �(��?@(/SO�FTPART/G�ENLINK?c�urrent=m�enupage,153,1���+��=�Oπ)��63=1�IE,2Pϣ�ȵ����*d�v�ed�it��PROG,A1��"�4�F���'��v�2����ߩ߻������ m��962 ��'�9�K�]������36�������p� ��
��.�@�R�d��������������� {�۱{�*<N` ru������� &8J\n� ������� "/4/F/X/j/|//�/ �/�/�/�/�/�/�/0? B?T?f?x?�??�?�? �?�?�?O��>OPO bOtO�O�O�?�O�O�O �O__�O:_L_^_p_ �_�_�_5_�_�_�_ o o$o�_HoZolo~o�o �o1o�o�o�o�o  2�oVhz��� ?���
��.�O +Od�v���������� ����*�<�ˏ`� r���������̟[�� ��&�8�J�ٟn��� ������ȯW����� "�4�F�X��|����� ��Ŀֿe�����0� B�T�?�Q��ϜϮ��� �������,�>�P� b���ߘߪ߼����� �߁��(�:�L�^�p� �ߔ���������}� ��$�6�H�Z�l�~�� �������������� �2DVhze����$UI_PANE�DATA 1L������  	�}/frh/gui��dev0.stm� M?conni�d=0 heig�ht=100&_�� ice=TP&�_lines=1�5&_colum�ns=4� fon�t=24&_pa�ge=whole�� �h�)pri9m/X  }[`����� )� ��#/
/G/Y/@/}/ d/�/�/�/�/�/�/?��/1?h��� �    �+��i�cgt?p/flex� ��?_width=(� �� 2�3� �1doub� 2;?8ual�?�?k O.O@OROdOvO?�O �O�O�O�O�O�O_*_ _N_5_r_Y_�_�_�_�_?= � �U�Oo $o6oHoZolo�_�oO �o�o�o�o�ouo2 D+hO���� ���
���@�'� d�v��_�_����Џ� ��Y�*��oN�`�r� ��������!�ޟş� �&�8��\�C����� y�����گ�ӯ��� ��F�X�j�|������ ĿֿI�����0�B� Tϻ�x�_ϜϮϕ��� �������,��P�b� I߆�mߪ��/���� ��(�:�L��p�� ����������U�� $��H�/�l�~�e��� ������������  DV���ߌ��� ��9
}�.@R dv����� �//�</#/`/r/ Y/�/}/�/�/�/�/c u&?8?J?\?n?�?�/ �?�?)�?�?�?O"O 4O�?XO?O|O�OuO�O �O�O�O�O_�O0_B_�)_f_M_�_�/?}���_�_�_�_
oo.o) �_So�5Boo�o�o�o �o�o@o�o�o! W>{b���� ����/��83;��$UI_POSTYPE  5�� 	 �;���a�QUICKMEN  p�����c�REST�ORE 1M5�  ��*defau�lt�;SIN�GLEԍPR�IMԏmwin�tpe,1,PROG,1<�p����� ��I���П����� ��<�N�`�r����"� �����ϯ��
��.� @��d�v�������O� п�����ï%�7� Iϻ��ϖϨϺ���o� ����&�8�J���n� �ߒߤ߶�a������� Y�"�4�F�X�j��� �������y����� 0�B�����a�s���� ����������,> Pbt��������SCRE��?���u1s]c�u2!3!U4!5!6!7!�8!�TATl��� ă5Y�USE1Rks#�U3�4�5�6��7�8�a�NDO_CFG Np���P�Qa�OP_CRM5  �U&a��PDd���None���_INFO 1O55f 0%��/ �8o/�/�/�/�/�/
? ?�/@?#?d?v?Y?�?�?�?�?��S!OFF?SET Rp�j!�?����!O3OEO WO�O{O�O�O�O�OO �O___J_A_S_�_ w_�_�_�Kŏ�]�_
o�
�_/o�8UFRA�M%�/P!RTOL_ABRTSoN#kb�ENBtoehGRP� 1S����Cz  A��c�a��o �o�o�o"v,>�cj��U�h#!�kMS�K  �ef!�kN6Pa%^)�%�_���e_EVNs`�t�&�v�2T�;
 }h#!UEVs`�!td:\ev�ent_user\�7�C7<�o� YFq�/�SP5�:��spotweldl�!C6��r���#�t!�K�	�>�� q��-��q���Q�c� ܟ�� �����ϟH�� l��)�_�����د�� ��˯ ��D���z� %�����[�m�濑�
����Ǻ�WRK 2U�a8�nπ� \ϥϷϒ������� �#���G�Y�4�}ߏ� j߳��ߠ���������1��B�g�y��$V�ARS_CONFuI�V�; FP�����CMR�b2�\�;xy� 	�$ ��01: S�C130EF2 Q*�	����X�ȸ�p�  #!?��p@pp"p�z� o]�g����@����������`�u�A����,�? B���G� K��l���_�� �����2� hSe�Q�����IA_WOF�]<^-˶,		�Q;%|/+'G�P �> ����RTWINU_RL ?�������/�/�/�/�/��/�SIONTM;OU� ��%��^S۳�S���@�a FR�:\�#\DATA�؏  �� wUD166LOGC?7  \9EXh?'q�' B@ ���2{1U��?{1�?��?θ � n?6  ������2�zt�`F��  =���BA��?@>|=TRAIN�?A4QB�d�CpBEFF�/B�0�(��_� (��I�M��O�O�O __P_>_t_b_|_�_��_�_�_�_�(_GE23`�/C�
�`'pX4b
g�0RE!0a�i\���LEXdb�����1-e�/VMPHASE  ����C ��RTD_�FILTER 2]c� �&��T� �o+=Oas �����o�������1�C�U�g��)S�HIFTMENU� 1d�K
 <b�<%�?ŏ2���� ɏ�ُ�8��!�n� E�W�}��������ß�՟"���	LIV�E/SNA��%?vsfliv�n4����# SETyU��W�menum��r��ѯ�"��3e�`+|�MO3ftn�-z��ZD�gQm˳�<�A�P�$WA�ITDINEND�8L!�k�OK  !�醼 :��S����wTIM5���Gr�͔�%˴��ӿx�򿆸RELE�a�5��k��/6m�_ACCTJ�4� !��_?17 h��%�5�<����RDIS��ο�$XVRna�itn�$ZABCv��1jQk ,�@r�2=��-ZIP2kQo���)����MPCF_G 1l��l!0L"��q�7�MP��m����P�������`��*�  ��f<�(G�3ޙ���?��6� 168Ÿ6�ff�H��C	���	(>�B��h��0�Q�����?����0B��r;T�ǯo@�S&������
�?�.�@�?�m�p9�������C���@�D"(>��N��a�3�]��2�� @l�PJ\r���D�)O�4%:��\�[(`68<_�6W�l����?�������0G�g8���Ea��'��J�p`n���_CYLIND��aoR� �p6? ,(  *o��w3l����  ��//'.iJ/�n/ U/g/�/��/�/�/// ?�/�/F?-?j?Q?�/��?�?�Cp*� �g��?L^���6O@!OZO?I�?�O?G��A�A�=SPHER/E 2qO�?�O T?�O_�O:_�?�Op_ �_�/�_E_+_�_�_ o �_Y_6oHo�_�_~o�_ �o�o�o�oo�o 6��ZZ�� ��