��   �A��*SYST�EM*��V9.1�035 7/1�9/2017 �A 	  ����PASSNAM�E_T   0� $+ �$'WORD  �? LEVEL � $TI- OU�TT��&F/�� $SET�UPJPROGR�AMJINSTA�LLJY  ?$CURR_O��USER�NUM��STSTOP_TPCHG V oLOG_P NT��N�  6 CO�UNT_DOWN��$ENB_P�CMPWD� $kDV_� IN� �$C� CRE���A RM9� T9DIAG9(�>LVCHK FULLM/�Y{XT�CNTDޏMENU�AU�TO+�FG_D�SP�RLS�U��BURYBAN��!eENC/�  CRY�PTE � ο��$$CL(  ? ���K!��� T @ V� ION�H(  ���\!IRTUA�� J/�$DCS_7COD?���O%��  W�'_S+  �*�� � �&��A91�"�!�	 
 $ R!�� =?"?0?F?T? j?x?�?�?�?�?�?�?��?OO,OBO���#S+UP� �*�DOVO�#FvO�O�O��  �L�A���_ � �� V�[t&��j���D�O^_��W_���t �V�U�YcELU�GH 1�) t �)�_�_ oo+o=oOoaoso�o �o�o�o�'�_�o�o 1CUgy�� ���o��	��-� ?�Q�c�u��������� �����)�;�M� _�q���������˟ڏ ���%�7�I�[�m� �������ǯ֟֯�� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛϭ� ���������+�=� O�a�s߅ߗߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1CUgy�� �����%