��   K�A��*SYST�EM*��V9.1�0185 12�/11/2019� A 	  ����CELL_�GRP_T  � � $'FR�AME $�MOUNT_LO�CCCF_MET�HOD  $�CPY_SRC_�IDX_PLATFRM_OFSC�tDIM_ $B�ASE{ FSET�C��AUX_O�RDER  � �XYZ_M�AP �� ~�LENGTH��TTCH_GP_�M~ a AUTOR�AIL_���$�$CLASS  ������D���DVERSI�ON � �i/IRT�UAL-9LO�OR G��DD3<x$?�������k,  1 <DwX< y�����C�����	/��Z�Zm//��/_/�/�/�/$ ��/�/	?';�$M�NU>A\"� � <�����3���g0��6 �7"!ik0�4x0s1�D�B� ��zP%$5{D-5!5�G.5!O�D*w1w0;�0�/s1º�+��?��Pv�95/ �?���?�?#O	O+OYO ?OqO�OuO�O�O�O�O��O_�O%_C_)_97N_UM  �����w92TOOLC?�\ 
Y;)/Y_"v�7_�_	o1_o?o %o7oYo�omo�o�o�o �o�o�o�o;!C qWy����� sV�Q�Vy�[