��   ��A��*SYST�EM*��V9.1�0185 12�/11/2019� A 
  ����DRYRU�N_T  4� $'ENB � $NUM_�PORTA ES�U@$STAT�E P TCOLu_��PMPMCm�GRP_MASK�ZE� OTION�NLOG_INF�ONiAVcFL�TR_EMPTY�d $PROD_�_ L �ESTOP�_DSBLAPOW_RECOVA�OPR�SAW_�� G %$I�NIT	RESUME_TYPEN�DIST_DIF}FA $ORN4 1� d =R��&J�_  4 u$(F3IDX��_ICI���MIX_BG-yy
_NAMc �MODc_US�d�IFY_TIv� �MKR-�  $LI�Nc   "_SIZc�� �. �X $USE_FLC 3!�8:&iF*SIMA7#�QC#QBn'SCAmN�AX�+IN�*}I��_COUNr�RO( ��!_TM�R_VA�g#h>�ia �'` �����1�+WA-R�$�H�!�#�N3CH�PEX�$O�!PR�'Iovq6�OoATH-� P $ENGABL+�0�BT��$$CL�ASS  �S���1��5��5�0�VERS��7  �iAIRTU� �?@'|/ 0E5���E����@kF1@�1pE��%�1�O���O��O����AEI2LK �O+_=_O_ a_s_�_�_�_�_�_�_ �_oo'o9o�O)W�?HW@ @��zj�0�o�o�i�� � 2LI G 4%Ho�o��mA }A�o+
Oa@� �v������ '���]�<�}A�c$"P+ �k�K@����pA��X��0A@�N �����0�B�T�f� x�����������pF}A Ձ}A����*�<�N� `�r���������̯ޯ��4hM��C� 2�lՏ;�M�_�q� ��������˿ݿ�� �Ԝ-�F�X�j�|ώ� �ϲ����������� )�B�T�f�xߊߜ߮� ����������,�7� P�b�t������� ������(�3�E�^� p���������������  $6A�Zl~ �������  2DOhz�� �����
//./ @/K]v/�/�/�/�/ �/�/�/??*?<?N? Qh�4�0���?=@