��   K�A��*SYST�EM*��V9.1�035 7/1�9/2017 �A 	  ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_���$$C�LASS  ������D��D�VERSION�  ���/IRTUA�L-9LOOR� G��DD<x$?������kn,  1 <DwX< y�����C�����	/��Z�Zm//�/_/p�/�/�/$ �/��/	?';�$MNU�>A\"�  <������3��g0��6 �"!�ik0�4x0s1D��B� ��zP%$5D-�5!5�G.5!�SD*w1w0;�0/s1�º�+���Pv�95/�?�� �?�?#O	O+OYO?OqO �OuO�O�O�O�O�O_��O%_C_)_97NUM  ����w92�TOOLC?\ y
Y;)-4��5�����PSQ,�Va�kBCv�7_ Y_	o1_o?o%o7oYo �omo�o�o�o�o�o�o �o;!CqWy �����sV�Q�V y�[