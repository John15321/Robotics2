��   v��A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����UI_CO�NFIG_T � x L$NU�M_MENUS � 9* NEC�TCRECOVE�R>CCOLOR�_CRR:EXT�STAT��$T{OP>_IDXC�MEM_LIMI�R$DBGLV�L�POPUP_�MASK�zA � $DUMMwY73�ODE�
]4CFOCA ��5CPS)C��\g HAN� � �TIMEOU�P�IPESIZE �� MWIN�P�ANEMAP� s � � FAVB ?� 
$HL�7_DIQ?� q�ELEMZ�URȩ l� Ss�$7HMI�RO+\�W ADONLY�� �TOUCH�PROOMM�O#?$�ALA�R< �FILVE9W�	ENB=�%%fC 1"USE�R:)FCTN:)W�I�� I* _E�D�l"V!_TIT�L� 1"COO�RDF<#LOCK�6%�$F%�!b"EBFOR�? �"e&1
�"�%�!BA�!j ���!BG�#�!hI{NSR$IO}�7PM�X_PK�T?$IHEL�P� ME�#BLN=KC=ENAB�!? �SIPMANUA�L4"="�BEE`Y?$�=&q!EDy#�M0IP0q!�JWqD�D7�DSB�V� GTB9I�:J�<wSTYf2$Iv!q_Gv!k FKE��FHTML�_wNAM�#DIMC4|:1]ABRIGH83s oDJ7CH92%!FE�L0T_DEVICzg1&USTO_@  t @;AR$@PIDD�B�C�D*PAG� ?�hA�B�ISCREVuEF���GN��@$FLAG�@���&�1  h� 	$PWD_A�CCES� MA�8��hS:1�%)$�LABE� $	Tz jHP�3�R�}	4SUSRVI >1  < `�Rp*�R��QPRI��m� t1�PTRI�P�"m�$$CL�ASP ����a��R��R `\ S�I�	g � �iaIRT�s1	o`'2 L1���L1���R	 K,��?���aF1`�b�d~a����c��y`� � �o��
 �� a�o�o1CU �oz����� c�
��.�@�R�� v���������Џ�q� ��*�<�N�`�� ������̟ޟm��� &�8�J�\�n������� ��ȯگ�{��"�4� F�X�j���������Ŀ�ֿ���`TPTX��ʊ�)��� s �Ƅ��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg���Ϩ�Ⱥ��υ�&a�s�pwd���+�=�O߄�s� �ߗߩ߻���\���� �'�9�K����߁��`����������a��`��b�b�� ($p�-����T�?�x���a�a��c���g���l��k
���Th�ah�h���h�	f����������`���`  q���f q��*h#h�Fd��g�Xc�B 1)hR �\ _�b �REG VE�D]���who�lemod.ht}m�	singl	�doub �trip8browsQ��� ��u���//�@/���dev�.sl�/3� 1�,	t�/_�/;/i/ ??/?�/S?e?w?�?�?�?� H`�?�?  OO$O6OHOZOlO~O�F @�?�O�O�O�O �O_�F�	�?�?;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo oM'�o�o�o�o�o�o +=Oas� ��������? >�P�b�t��������� Ώ���O�����L� ^�_'_�������ş �����6�1�C�U� ~�y�����Ư��ӯ�o ���-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�-��Ϭ� ����������*�<� 7�`�r�A�Sߨߺ�q� ��i�����!�J�E� W�i��������� ����"��/���O�I� w��������������� +=Oas� ������, >Pbt���߼ ���//����� ^/Y/k/}/�/�/�/�/ �/�/�/?6?1?C?U? ~?y?�?Y��?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _�R_d_v_�_�_�_ �_�_�_�_�o*o�_�o`oro�j�$UI�_TOPMENU� 1K`�aR 
d�a�*Q)*defa�ult5_]*�level0 * [	 �o�0��o'rtpio�[23]�8tpst[1[x)w9��o	�=h58E�01_l.png���6menu5�y�p�13�z��zb	�4���q��]� ��������̏ޏ)Rr����+�=�O�a����prim=�pa�ge,1422,1h�����şן����1�C�U�g����|�class,5�p�����ɯۯ�����13��*�<�N�`�4r���|�53�������ҿ�����|�8 ��1�C�U�g�y�����@����������"Y�` �a�o/��m!ηq�Y��w�avtyl}Tfqm�f[0nl�	��c�[164[w��59@[x�qG���/��29� �o�%�1���{��m� �!�����0�B��� f�x���������O������,>����2 P�����\�� '9K�������������1���/$/6/H/Z/��~|�ainedi'���/�/�/�/�/��c�onfig=si�ngle&|�wintp���/$?6?H? Z?!Z�a�h?�?�e�? �;��?�?�?OO+O =OOO�?[O�O�O�O�O �O�O�O_a�%_L_^_ p_�_�_�_���_�_�_  oo$o�_HoZolo~o �o�o1o�o�o�o�o  2�oVhz�� �?���
��.� �@�d�v��������� M�����*�<�ˏ�`�r���������^ ��;�M�sc�_;����s��X�}���e�u ��0���P��t���4�j�X�6e�u7 �����ｿϿ��� P�)�;�M�_�qσ�� �Ϲ����������"�1�M�_�q߃� �ߠϹ��������� ��7�I�[�m���� ����������!�����6(�]�o��������$��74�������)t<ϯ\�5	TPTX[209©|Dw24§J����w18����
�02��A#��[�tv`�RdvL0�K1���5S�:�$treevi�ew3��3��&d�ual=o'81,26,4�O/a/ s/2�/�/�/�/�/�/ �/?'?9?K?]?o?��;/��53$/6$�� �?�?�?
?#O5OGOYO kO}OO�O�O�O�O�O��O�?�?��1�?6$2p�f_x_�_ �6_��edit��>_P_ �_�_o��/���_�S ooo�o�oB�o�o� �oA�o�+= Oas��o��� ����(�9���Q� x���������ҏ�O�� ��,�>�P�ߏt��� ������Ο]����� (�:�L�^�ퟂ����� ��ʯܯk� ��$�6� H�Z��l�������ƿ ؿ�y�� �2�D�V� h����Ϟϰ������� �o�o��o@ߧE�c� u߇ߙ߽߬�����O� ���)�<�M�_�q�� ��W���������&� 8���\�n��������� E�������"4�� Xj|����S ��0B�f x����O�� //,/>/P/�t/�/ �/�/�/�/]/�/?? (?:?L?��߂?1ߦ? ���?�?�?�?O$O 5OGO�?SO}O�O�O�O �O�O�O�O��2_D_V_ h_z_�_�_�/�_�_�_ �_
oo�_@oRodovo �o�o)o�o�o�o�o *�oN`r�� �7�����&� �J�\�n��������� E�ڏ����"�4�Ï X�j�|�������a?s? 蟗?�sO_/�A�S� e�w����������� ����,�=�O�a�#_ ������ο��=�� (�:�L�^�pς�Ϧ� �������� ߏ�$�6� H�Z�l�~�ߐߴ��� ��������2�D�V� h�z���������� ��
����@�R�d�v� ����)����������ƚԔ*def�ault%��*?level8�ٯ�w���? t?pst[1]�	��y�tpio[#23���u����J\menu7_l.png_M|13��5�h{�y4�u6� ��//'/9/K/]/�� �/�/�/�/�/�/j/�/�?#?5?G?Y?k?�"�prim=|page,74,1p?@�?�?�?�?�?�"�6�class,13 �?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo�]ooo�o`�$UI�_USERVIE�W 1֑֑�R 
�A��o��o�o[m�o '9K] �� ���l���#� 5��oB�T�f������ ŏ׏鏌���1�C� U�g�
���������ӟ ~�����v�?�Q�c� u���*�����ϯ�� ���)�;�M�_�
�� ~������ݿ��� %�ȿI�[�m�ϑ�4� ���������Ϩ�
�� .ߠ�i�{ߍߟ߱�T� ��������/���S� e�w���Fߨ���� >���+�=�O���s� ��������^����� '����FX��| ������# 5GY�}��� �p���h1/C/ U/g/y//�/�/�/�/ �/�/�/?-???Q?c? /p?�?�??�?�?�? OO�?;OMO_OqO�O &O�O�O�O�O�O�?�O _ _�OD_m__�_�_ �_X_�_�_�_o!o�_ EoWoio{o�o0h