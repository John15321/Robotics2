��   ��A��*SYST�EM*��V9.1�035 7/1�9/2017 �A 
  ����DRYRUN_�T  4 �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	RESUME�_TYPENDIST_DIFFA $ORN41� 8d =R��&J�_  4 u$(F3IDX��_ICI  �MIX_BG-yy
_NAMc �MODc_US�d�IFY_TI�� ��MKR�-  $L{INc   "_SIZcg�� ��. X $?USE_FLC �3!�:&iF*SIM�A7#QC#QBn'S�CAN�AX�+I�N�*I��_COU�NrRO( ��!_?TMR_VA�g#h>�ia  �'` ����1�+�WAR�$�H4�!�#N3CH�cPE�$O�!PR�'�Ioq6�OoAT�H- P $ENABL+��0BTf�$$�CLASS  O����1��5��=5�0VERS��7�  �=�AIRTU� �?�@'/ 0E5�������@kF!1@�1pE��%�1�O���O�O����AEI;2LK �O+_ =_O_a_s_�_�_�_�_ �_�_�_oo'o9o�O�)W?HW@ ��zj�0�o�o�i��� � 2LI  4%Ho�o��mA}A�o+
Oa @��v���� ��'���]�<�}A@�c$"+ �k�K@��1��pA��XyA0A @�N�����0�B� T�f�x����������� pF}AՁ}A����*� <�N�`�r����������̯ޯ�4hM��C� 2Ђ�hՏ;�M� _�q���������˿ݿ ���Ԝ-�F�X�j� |ώϠϲ��������� ��)�B�T�f�xߊ� �߮����������� ,�7�P�b�t���� ����������(�3� E�^�p����������� ���� $6A�Z l~������ � 2DOhz �������
/ /./@/K]v/�/�/ �/�/�/�/�/??*? <?N?Qh�4�0���?=@