��   ��A��*SYST�EM*��V9.1�035 7/1�9/2017 �A 
  ����DRYRUN_�T  4 �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	RESUME�_TYPENDIST_DIFFA $ORN41� 8d =R��&J�_  4 u$(F3IDX�̈_ICIfMI/X_BG-y
�_NAMc MO�Dc_USd�I�FY_TI� �MKR- � $LINc  � "_SIZ�c�� �. X� $USE_FLC 3!�:&iF*SIMA7#QC#Q�Bn'SCAN�A�X�+IN�*I��_oCOUNrRO( ���!_TMR_V1A�g#h> �ia �'` �����1�+WAR��$�H�!�#N3CH�PE�$O�!�PR�'Ioq6�O�oATH- P� $ENABL+�0BTf��$$CLASS  ����1���5��5�0VER�S��7 � ��AIRT�U� �?@'/ 0E�5�������@kF1@�1pE���%�1�O���O�O�����AEI2LK �O+_=_O_a_s_�_ �_�_�_�_�_�_oo`'o9o�O)W?HW@ ��zj�0Ȋo�o�i�� � 2�LI  4%Ho�o��mA}A�o+ 
Oa@��v� �����'��� ]�<�}A�c$"+ �k�K�@����pA��XmA0A@�N���� �0�B�T�f�x����� ������pF}AՁ}A�� ��*�<�N�`�r����������̯ޯ�4hM���C� 2�l Տ;�M�_�q������� ��˿ݿ���Ԝ-� F�X�j�|ώϠϲ��� ��������)�B�T� f�xߊߜ߮������� ����,�7�P�b�t� ������������ �(�3�E�^�p����� ���������� $ 6A�Zl~��� ���� 2D Ohz����� ��
//./@/K] v/�/�/�/�/�/�/�/ ??*?<?N?Qh�4�0 ���?=@