��   �A��*SYST�EM*��V9.1�0185 12�/11/2019� A   ����BIN_C�FG_T   �X 	$ENTR�IES  $�Q0FP?NG1�F1O2F2OP�z ?CNETG����DHCP_C�TRL.  0{ 7 ABLE? �$IPUS�R�ETRAT�$SETHOST��NSS* 8��D�FACE_�NUM? $DBG_LEVEL��OM_NAM� �!� FT� =@� LOG_8	,�CMO>$DN�LD_FILTE�R�SUBDIRCAPC��8 .� 4� H{A�DDRTYP�H NGTH��� �z +LSq� D $ROB�OTIG �PEEyR�� MASK��MRU~OMGD�EV��PINF�O�  $�$$TI ���RCM+T A$( /�QSIZ�!S� �TATUS_%$�MAILSERV~ $PLAN� �<$LIN<�$CLU��<${TO�P$CC�&sFR�&YJEC|!}Z%ENB � �ALAR:!B�TQP,�#,V8 S��_$VAR�)M��ON�&���&APPL�&PA� �%��''POR�Y#_�!�"�ALERT�&i2U�RL }Z3A�TTAC��0ER�R_THROU3UaS�9H!�8� CH- �c%�4MAX?WS�_|1��1MO	D��1I�  �1o �(�1PWD  Ɵ LA��0�ND��1TRYFDEL�A-C�0G'AERS�I��1Q'ROBIC�LK_HM 0Q'� X�ML+ 3SGFReMU3T� !OUU3f G_�-COP1�F33�AQ'C[2�%�B_AU�� 9 R�!�UPDb&PCO�U{!�CFO 2 
$V*W�@�c%ACC_HYQSN}A�UMMY1oW�2"$DM* �$DIS��SN,#	3 �	o!�"�%"_WI�CTZ�_INDE�3�PO�FF� ~UR�YD���S�  
 �t Z!RT�0N�(cD�)bHOUU#E%A/fVa>fVaMf�LOCA� #$�NS0H_HE����@I�/  dκPARPH&�_IPF�W_* O�F�PQFAsD90��VHO_� 5R42PyS�a?�TEL�G P����90WORAXQE�� LVO#�FS1��ICE�[p� ��$�c  ��)�zq��
��
op�PyS�Axw# k�i�qIz0ALw��q'0 �x
���F������p�r�u�]$� 2�{ ���r#���� �}��!�qi����$� _?FLTR  �y�pW �������!�}�$�}2}��boSHAR� 1�yE Pe���t
� G�6�k�.���R���v� ������П1���U� �y�<���`�r�ӯ�� �����ޯ?���u� 8���\�����ῤ�ڿ ��;���_�"σ�F� ��jϸ��Ϡ����%� ��I��m�0�Bߣ�f� �ߊ��߮������E� �i�,��P��t���������/���z _�LUA1��x!�1.j�08���i�1|z���255.��Lq�����uh�2o���������������3 ����^ 1C��4_��� ������5���N�!3��6O���u�ș����QJ��a��a� ��(�� OQ� '��<a/ �/�/{/�/�/�/�/?&?��P?V?h?z?9? �?�?�?�?�?�?
OO���?���ufOQL�
ZDT Status�?uO�O�O�O���}iRCon�nect: ir�c�D//alert�N&_8_J_\_�G�O��_�_�_�_�_�_��r�sP 2ـd���_ o1oCoUogoyo�o�o��o�o�o�o�o�s$$�c962b37a�-1ac0-eb�2a-f1c7-�8c6eb5f01a8c  (y_�J�On������ـP(�X"�rZJ��u3 �v[C] )�,$ e"�ـ[��M�4�q� X�~�����ˏ���� �%��I�0�B��f�h�������w�W�n8 DM_=!W��G�SNTP�	��%��-����������K�4#��USTOM 
�2F��W  �3$_TCPIP��aXHO%S"��ELO��W�T!�E�H!�Tb���rj_3_tpdQO \�~�!KCL��������v!CR�TY�G���O"(�!�CONS�� ���ib_smon����